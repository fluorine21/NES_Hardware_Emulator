

package vram_listing;


integer spram_listing[64] = 
{
//Sprite 0
8'h00, 8'h00, //row 0
8'h01, 8'h00, // Tile 1F
8'h02, 8'h00, // Attribute bytes
8'h03, 8'h00, //Col 0

//Sprite 1
8'h04, 8'h08, //row 0
8'h05, 8'h00, // Tile 1F
8'h06, 8'h01, // Attribute bytes
8'h07, 8'h08, //Col 8

//Sprite 2
8'h08, 8'h10, //row 0
8'h09, 8'h00, // Tile 1F
8'h0A, 8'h02, // Attribute bytes
8'h0B, 8'h10, //Col 16

//Sprite 3
8'h0C, 8'h18, //row 0
8'h0D, 8'h00, // Tile 1F
8'h0E, 8'h03, // Attribute bytes
8'h0F, 8'h18, //Col 24

//Sprite 4
8'h10, 8'h20, //row 0
8'h11, 8'h00, // Tile 1F
8'h12, 8'h00, // Attribute bytes
8'h13, 8'h20, //Col 32

//Sprite 5
8'h14, 8'h28, //row 0
8'h15, 8'h00, // Tile 1F
8'h16, 8'h01, // Attribute bytes
8'h17, 8'h28, //Col 40

//Sprite 6
8'h18, 8'h30, //row 0
8'h19, 8'h00, // Tile 1F
8'h1A, 8'h02, // Attribute bytes
8'h1B, 8'h30, //Col 48

//Sprite 7
8'h1C, 8'h38, //row 0
8'h1D, 8'h00, // Tile 1F
8'h1E, 8'h03, // Attribute bytes
8'h1F, 8'h38 //Col 56
};



integer vram_listing[] = 
{


16'h0000, 16'hFFFF,
16'h0001, 16'hFFFF,
16'h0002, 16'hFFFF,
16'h0003, 16'hFFFF,
16'h0004, 16'hFFFF,
16'h0005, 16'hFFFF,
16'h0006, 16'hFFFF,
16'h0007, 16'hFFFF,
16'h0008, 16'hFFFF,
16'h0009, 16'hFFFF,
16'h000A, 16'hFFFF,
16'h000B, 16'hFFFF,
16'h000C, 16'hFFFF,
16'h000D, 16'hFFFF,
16'h000E, 16'hFFFF,
16'h000F, 16'hFFFF,
16'h0010, 16'hFFFF,
16'h0011, 16'hFFFF,
16'h0012, 16'hFFFF,
16'h0013, 16'hFFFF,
16'h0014, 16'hFFFF,
16'h0015, 16'hFFFF,
16'h0016, 16'hFFFF,
16'h0017, 16'hFFFF,
16'h0018, 16'hFFFF,
16'h0019, 16'hFFFF,
16'h001A, 16'hFFFF,
16'h001B, 16'hFFFF,
16'h001C, 16'hFFFF,
16'h001D, 16'hFFFF,
16'h001E, 16'hFFFF,
16'h001F, 16'hFFFF,
16'h0020, 16'hFFFF,
16'h0021, 16'hFFFF,
16'h0022, 16'hFFFF,
16'h0023, 16'hFFFF,
16'h0024, 16'hFFFF,
16'h0025, 16'hFFFF,
16'h0026, 16'hFFFF,
16'h0027, 16'hFFFF,
16'h0028, 16'hFFFF,
16'h0029, 16'hFFFF,
16'h002A, 16'hFFFF,
16'h002B, 16'hFFFF,
16'h002C, 16'hFFFF,
16'h002D, 16'hFFFF,
16'h002E, 16'hFFFF,
16'h002F, 16'hFFFF,
16'h0030, 16'hFFFF,
16'h0031, 16'hFFFF,
16'h0032, 16'hFFFF,
16'h0033, 16'hFFFF,
16'h0034, 16'hFFFF,
16'h0035, 16'hFFFF,
16'h0036, 16'hFFFF,
16'h0037, 16'hFFFF,
16'h0038, 16'hFFFF,
16'h0039, 16'hFFFF,
16'h003A, 16'hFFFF,
16'h003B, 16'hFFFF,
16'h003C, 16'hFFFF,
16'h003D, 16'hFFFF,
16'h003E, 16'hFFFF,
16'h003F, 16'hFFFF,
16'h0040, 16'hFFFF,
16'h0041, 16'hFFFF,
16'h0042, 16'hFFFF,
16'h0043, 16'hFFFF,
16'h0044, 16'hFFFF,
16'h0045, 16'hFFFF,
16'h0046, 16'hFFFF,
16'h0047, 16'hFFFF,
16'h0048, 16'hFFFF,
16'h0049, 16'hFFFF,
16'h004A, 16'hFFFF,
16'h004B, 16'hFFFF,
16'h004C, 16'hFFFF,
16'h004D, 16'hFFFF,
16'h004E, 16'hFFFF,
16'h004F, 16'hFFFF,
16'h0050, 16'hFFFF,
16'h0051, 16'hFFFF,
16'h0052, 16'hFFFF,
16'h0053, 16'hFFFF,
16'h0054, 16'hFFFF,
16'h0055, 16'hFFFF,
16'h0056, 16'hFFFF,
16'h0057, 16'hFFFF,
16'h0058, 16'hFFFF,
16'h0059, 16'hFFFF,
16'h005A, 16'hFFFF,
16'h005B, 16'hFFFF,
16'h005C, 16'hFFFF,
16'h005D, 16'hFFFF,
16'h005E, 16'hFFFF,
16'h005F, 16'hFFFF,
16'h0060, 16'hFFFF,
16'h0061, 16'hFFFF,
16'h0062, 16'hFFFF,
16'h0063, 16'hFFFF,
16'h0064, 16'hFFFF,
16'h0065, 16'hFFFF,
16'h0066, 16'hFFFF,
16'h0067, 16'hFFFF,
16'h0068, 16'hFFFF,
16'h0069, 16'hFFFF,
16'h006A, 16'hFFFF,
16'h006B, 16'hFFFF,
16'h006C, 16'hFFFF,
16'h006D, 16'hFFFF,
16'h006E, 16'hFFFF,
16'h006F, 16'hFFFF,
16'h0070, 16'hFFFF,
16'h0071, 16'hFFFF,
16'h0072, 16'hFFFF,
16'h0073, 16'hFFFF,
16'h0074, 16'hFFFF,
16'h0075, 16'hFFFF,
16'h0076, 16'hFFFF,
16'h0077, 16'hFFFF,
16'h0078, 16'hFFFF,
16'h0079, 16'hFFFF,
16'h007A, 16'hFFFF,
16'h007B, 16'hFFFF,
16'h007C, 16'hFFFF,
16'h007D, 16'hFFFF,
16'h007E, 16'hFFFF,
16'h007F, 16'hFFFF,
16'h0080, 16'hFFFF,
16'h0081, 16'hFFFF,
16'h0082, 16'hFFFF,
16'h0083, 16'hFFFF,
16'h0084, 16'hFFFF,
16'h0085, 16'hFFFF,
16'h0086, 16'hFFFF,
16'h0087, 16'hFFFF,
16'h0088, 16'hFFFF,
16'h0089, 16'hFFFF,
16'h008A, 16'hFFFF,
16'h008B, 16'hFFFF,
16'h008C, 16'hFFFF,
16'h008D, 16'hFFFF,
16'h008E, 16'hFFFF,
16'h008F, 16'hFFFF,
16'h0090, 16'hFFFF,
16'h0091, 16'hFFFF,
16'h0092, 16'hFFFF,
16'h0093, 16'hFFFF,
16'h0094, 16'hFFFF,
16'h0095, 16'hFFFF,
16'h0096, 16'hFFFF,
16'h0097, 16'hFFFF,
16'h0098, 16'hFFFF,
16'h0099, 16'hFFFF,
16'h009A, 16'hFFFF,
16'h009B, 16'hFFFF,
16'h009C, 16'hFFFF,
16'h009D, 16'hFFFF,
16'h009E, 16'hFFFF,
16'h009F, 16'hFFFF,
16'h00A0, 16'hFFFF,
16'h00A1, 16'hFFFF,
16'h00A2, 16'hFFFF,
16'h00A3, 16'hFFFF,
16'h00A4, 16'hFFFF,
16'h00A5, 16'hFFFF,
16'h00A6, 16'hFFFF,
16'h00A7, 16'hFFFF,
16'h00A8, 16'hFFFF,
16'h00A9, 16'hFFFF,
16'h00AA, 16'hFFFF,
16'h00AB, 16'hFFFF,
16'h00AC, 16'hFFFF,
16'h00AD, 16'hFFFF,
16'h00AE, 16'hFFFF,
16'h00AF, 16'hFFFF,
16'h00B0, 16'hFFFF,
16'h00B1, 16'hFFFF,
16'h00B2, 16'hFFFF,
16'h00B3, 16'hFFFF,
16'h00B4, 16'hFFFF,
16'h00B5, 16'hFFFF,
16'h00B6, 16'hFFFF,
16'h00B7, 16'hFFFF,
16'h00B8, 16'hFFFF,
16'h00B9, 16'hFFFF,
16'h00BA, 16'hFFFF,
16'h00BB, 16'hFFFF,
16'h00BC, 16'hFFFF,
16'h00BD, 16'hFFFF,
16'h00BE, 16'hFFFF,
16'h00BF, 16'hFFFF,
16'h00C0, 16'hFFFF,
16'h00C1, 16'hFFFF,
16'h00C2, 16'hFFFF,
16'h00C3, 16'hFFFF,
16'h00C4, 16'hFFFF,
16'h00C5, 16'hFFFF,
16'h00C6, 16'hFFFF,
16'h00C7, 16'hFFFF,
16'h00C8, 16'hFFFF,
16'h00C9, 16'hFFFF,
16'h00CA, 16'hFFFF,
16'h00CB, 16'hFFFF,
16'h00CC, 16'hFFFF,
16'h00CD, 16'hFFFF,
16'h00CE, 16'hFFFF,
16'h00CF, 16'hFFFF,
16'h00D0, 16'hFFFF,
16'h00D1, 16'hFFFF,
16'h00D2, 16'hFFFF,
16'h00D3, 16'hFFFF,
16'h00D4, 16'hFFFF,
16'h00D5, 16'hFFFF,
16'h00D6, 16'hFFFF,
16'h00D7, 16'hFFFF,
16'h00D8, 16'hFFFF,
16'h00D9, 16'hFFFF,
16'h00DA, 16'hFFFF,
16'h00DB, 16'hFFFF,
16'h00DC, 16'hFFFF,
16'h00DD, 16'hFFFF,
16'h00DE, 16'hFFFF,
16'h00DF, 16'hFFFF,
16'h00E0, 16'hFFFF,
16'h00E1, 16'hFFFF,
16'h00E2, 16'hFFFF,
16'h00E3, 16'hFFFF,
16'h00E4, 16'hFFFF,
16'h00E5, 16'hFFFF,
16'h00E6, 16'hFFFF,
16'h00E7, 16'hFFFF,
16'h00E8, 16'hFFFF,
16'h00E9, 16'hFFFF,
16'h00EA, 16'hFFFF,
16'h00EB, 16'hFFFF,
16'h00EC, 16'hFFFF,
16'h00ED, 16'hFFFF,
16'h00EE, 16'hFFFF,
16'h00EF, 16'hFFFF,
16'h00F0, 16'hFFFF,
16'h00F1, 16'hFFFF,
16'h00F2, 16'hFFFF,
16'h00F3, 16'hFFFF,
16'h00F4, 16'hFFFF,
16'h00F5, 16'hFFFF,
16'h00F6, 16'hFFFF,
16'h00F7, 16'hFFFF,
16'h00F8, 16'hFFFF,
16'h00F9, 16'hFFFF,
16'h00FA, 16'hFFFF,
16'h00FB, 16'hFFFF,
16'h00FC, 16'hFFFF,
16'h00FD, 16'hFFFF,
16'h00FE, 16'hFFFF,
16'h00FF, 16'hFFFF,
16'h0100, 16'hFFFF,
16'h0101, 16'hFFFF,
16'h0102, 16'hFFFF,
16'h0103, 16'hFFFF,
16'h0104, 16'hFFFF,
16'h0105, 16'hFFFF,
16'h0106, 16'hFFFF,
16'h0107, 16'hFFFF,
16'h0108, 16'hFFFF,
16'h0109, 16'hFFFF,
16'h010A, 16'hFFFF,
16'h010B, 16'hFFFF,
16'h010C, 16'hFFFF,
16'h010D, 16'hFFFF,
16'h010E, 16'hFFFF,
16'h010F, 16'hFFFF,
16'h0110, 16'hFFFF,
16'h0111, 16'hFFFF,
16'h0112, 16'hFFFF,
16'h0113, 16'hFFFF,
16'h0114, 16'hFFFF,
16'h0115, 16'hFFFF,
16'h0116, 16'hFFFF,
16'h0117, 16'hFFFF,
16'h0118, 16'hFFFF,
16'h0119, 16'hFFFF,
16'h011A, 16'hFFFF,
16'h011B, 16'hFFFF,
16'h011C, 16'hFFFF,
16'h011D, 16'hFFFF,
16'h011E, 16'hFFFF,
16'h011F, 16'hFFFF,
16'h0120, 16'hFFFF,
16'h0121, 16'hFFFF,
16'h0122, 16'hFFFF,
16'h0123, 16'hFFFF,
16'h0124, 16'hFFFF,
16'h0125, 16'hFFFF,
16'h0126, 16'hFFFF,
16'h0127, 16'hFFFF,
16'h0128, 16'hFFFF,
16'h0129, 16'hFFFF,
16'h012A, 16'hFFFF,
16'h012B, 16'hFFFF,
16'h012C, 16'hFFFF,
16'h012D, 16'hFFFF,
16'h012E, 16'hFFFF,
16'h012F, 16'hFFFF,
16'h0130, 16'hFFFF,
16'h0131, 16'hFFFF,
16'h0132, 16'hFFFF,
16'h0133, 16'hFFFF,
16'h0134, 16'hFFFF,
16'h0135, 16'hFFFF,
16'h0136, 16'hFFFF,
16'h0137, 16'hFFFF,
16'h0138, 16'hFFFF,
16'h0139, 16'hFFFF,
16'h013A, 16'hFFFF,
16'h013B, 16'hFFFF,
16'h013C, 16'hFFFF,
16'h013D, 16'hFFFF,
16'h013E, 16'hFFFF,
16'h013F, 16'hFFFF,
16'h0140, 16'hFFFF,
16'h0141, 16'hFFFF,
16'h0142, 16'hFFFF,
16'h0143, 16'hFFFF,
16'h0144, 16'hFFFF,
16'h0145, 16'hFFFF,
16'h0146, 16'hFFFF,
16'h0147, 16'hFFFF,
16'h0148, 16'hFFFF,
16'h0149, 16'hFFFF,
16'h014A, 16'hFFFF,
16'h014B, 16'hFFFF,
16'h014C, 16'hFFFF,
16'h014D, 16'hFFFF,
16'h014E, 16'hFFFF,
16'h014F, 16'hFFFF,
16'h0150, 16'hFFFF,
16'h0151, 16'hFFFF,
16'h0152, 16'hFFFF,
16'h0153, 16'hFFFF,
16'h0154, 16'hFFFF,
16'h0155, 16'hFFFF,
16'h0156, 16'hFFFF,
16'h0157, 16'hFFFF,
16'h0158, 16'hFFFF,
16'h0159, 16'hFFFF,
16'h015A, 16'hFFFF,
16'h015B, 16'hFFFF,
16'h015C, 16'hFFFF,
16'h015D, 16'hFFFF,
16'h015E, 16'hFFFF,
16'h015F, 16'hFFFF,
16'h0160, 16'hFFFF,
16'h0161, 16'hFFFF,
16'h0162, 16'hFFFF,
16'h0163, 16'hFFFF,
16'h0164, 16'hFFFF,
16'h0165, 16'hFFFF,
16'h0166, 16'hFFFF,
16'h0167, 16'hFFFF,
16'h0168, 16'hFFFF,
16'h0169, 16'hFFFF,
16'h016A, 16'hFFFF,
16'h016B, 16'hFFFF,
16'h016C, 16'hFFFF,
16'h016D, 16'hFFFF,
16'h016E, 16'hFFFF,
16'h016F, 16'hFFFF,
16'h0170, 16'hFFFF,
16'h0171, 16'hFFFF,
16'h0172, 16'hFFFF,
16'h0173, 16'hFFFF,
16'h0174, 16'hFFFF,
16'h0175, 16'hFFFF,
16'h0176, 16'hFFFF,
16'h0177, 16'hFFFF,
16'h0178, 16'hFFFF,
16'h0179, 16'hFFFF,
16'h017A, 16'hFFFF,
16'h017B, 16'hFFFF,
16'h017C, 16'hFFFF,
16'h017D, 16'hFFFF,
16'h017E, 16'hFFFF,
16'h017F, 16'hFFFF,
16'h0180, 16'hFFFF,
16'h0181, 16'hFFFF,
16'h0182, 16'hFFFF,
16'h0183, 16'hFFFF,
16'h0184, 16'hFFFF,
16'h0185, 16'hFFFF,
16'h0186, 16'hFFFF,
16'h0187, 16'hFFFF,
16'h0188, 16'hFFFF,
16'h0189, 16'hFFFF,
16'h018A, 16'hFFFF,
16'h018B, 16'hFFFF,
16'h018C, 16'hFFFF,
16'h018D, 16'hFFFF,
16'h018E, 16'hFFFF,
16'h018F, 16'hFFFF,
16'h0190, 16'hFFFF,
16'h0191, 16'hFFFF,
16'h0192, 16'hFFFF,
16'h0193, 16'hFFFF,
16'h0194, 16'hFFFF,
16'h0195, 16'hFFFF,
16'h0196, 16'hFFFF,
16'h0197, 16'hFFFF,
16'h0198, 16'hFFFF,
16'h0199, 16'hFFFF,
16'h019A, 16'hFFFF,
16'h019B, 16'hFFFF,
16'h019C, 16'hFFFF,
16'h019D, 16'hFFFF,
16'h019E, 16'hFFFF,
16'h019F, 16'hFFFF,
16'h01A0, 16'hFFFF,
16'h01A1, 16'hFFFF,
16'h01A2, 16'hFFFF,
16'h01A3, 16'hFFFF,
16'h01A4, 16'hFFFF,
16'h01A5, 16'hFFFF,
16'h01A6, 16'hFFFF,
16'h01A7, 16'hFFFF,
16'h01A8, 16'hFFFF,
16'h01A9, 16'hFFFF,
16'h01AA, 16'hFFFF,
16'h01AB, 16'hFFFF,
16'h01AC, 16'hFFFF,
16'h01AD, 16'hFFFF,
16'h01AE, 16'hFFFF,
16'h01AF, 16'hFFFF,
16'h01B0, 16'hFFFF,
16'h01B1, 16'hFFFF,
16'h01B2, 16'hFFFF,
16'h01B3, 16'hFFFF,
16'h01B4, 16'hFFFF,
16'h01B5, 16'hFFFF,
16'h01B6, 16'hFFFF,
16'h01B7, 16'hFFFF,
16'h01B8, 16'hFFFF,
16'h01B9, 16'hFFFF,
16'h01BA, 16'hFFFF,
16'h01BB, 16'hFFFF,
16'h01BC, 16'hFFFF,
16'h01BD, 16'hFFFF,
16'h01BE, 16'hFFFF,
16'h01BF, 16'hFFFF,
16'h01C0, 16'hFFFF,
16'h01C1, 16'hFFFF,
16'h01C2, 16'hFFFF,
16'h01C3, 16'hFFFF,
16'h01C4, 16'hFFFF,
16'h01C5, 16'hFFFF,
16'h01C6, 16'hFFFF,
16'h01C7, 16'hFFFF,
16'h01C8, 16'hFFFF,
16'h01C9, 16'hFFFF,
16'h01CA, 16'hFFFF,
16'h01CB, 16'hFFFF,
16'h01CC, 16'hFFFF,
16'h01CD, 16'hFFFF,
16'h01CE, 16'hFFFF,
16'h01CF, 16'hFFFF,
16'h01D0, 16'hFFFF,
16'h01D1, 16'hFFFF,
16'h01D2, 16'hFFFF,
16'h01D3, 16'hFFFF,
16'h01D4, 16'hFFFF,
16'h01D5, 16'hFFFF,
16'h01D6, 16'hFFFF,
16'h01D7, 16'hFFFF,
16'h01D8, 16'hFFFF,
16'h01D9, 16'hFFFF,
16'h01DA, 16'hFFFF,
16'h01DB, 16'hFFFF,
16'h01DC, 16'hFFFF,
16'h01DD, 16'hFFFF,
16'h01DE, 16'hFFFF,
16'h01DF, 16'hFFFF,
16'h01E0, 16'hFFFF,
16'h01E1, 16'hFFFF,
16'h01E2, 16'hFFFF,
16'h01E3, 16'hFFFF,
16'h01E4, 16'hFFFF,
16'h01E5, 16'hFFFF,
16'h01E6, 16'hFFFF,
16'h01E7, 16'hFFFF,
16'h01E8, 16'hFFFF,
16'h01E9, 16'hFFFF,
16'h01EA, 16'hFFFF,
16'h01EB, 16'hFFFF,
16'h01EC, 16'hFFFF,
16'h01ED, 16'hFFFF,
16'h01EE, 16'hFFFF,
16'h01EF, 16'hFFFF,
16'h01F0, 16'hFFFF,
16'h01F1, 16'hFFFF,
16'h01F2, 16'hFFFF,
16'h01F3, 16'hFFFF,
16'h01F4, 16'hFFFF,
16'h01F5, 16'hFFFF,
16'h01F6, 16'hFFFF,
16'h01F7, 16'hFFFF,
16'h01F8, 16'hFFFF,
16'h01F9, 16'hFFFF,
16'h01FA, 16'hFFFF,
16'h01FB, 16'hFFFF,
16'h01FC, 16'hFFFF,
16'h01FD, 16'hFFFF,
16'h01FE, 16'hFFFF,
16'h01FF, 16'hFFFF,
16'h0200, 16'hFFFF,
16'h0201, 16'hFFFF,
16'h0202, 16'hFFFF,
16'h0203, 16'hFFFF,
16'h0204, 16'hFFFF,
16'h0205, 16'hFFFF,
16'h0206, 16'hFFFF,
16'h0207, 16'hFFFF,
16'h0208, 16'hFFFF,
16'h0209, 16'hFFFF,
16'h020A, 16'hFFFF,
16'h020B, 16'hFFFF,
16'h020C, 16'hFFFF,
16'h020D, 16'hFFFF,
16'h020E, 16'hFFFF,
16'h020F, 16'hFFFF,
16'h0210, 16'hFFFF,
16'h0211, 16'hFFFF,
16'h0212, 16'hFFFF,
16'h0213, 16'hFFFF,
16'h0214, 16'hFFFF,
16'h0215, 16'hFFFF,
16'h0216, 16'hFFFF,
16'h0217, 16'hFFFF,
16'h0218, 16'hFFFF,
16'h0219, 16'hFFFF,
16'h021A, 16'hFFFF,
16'h021B, 16'hFFFF,
16'h021C, 16'hFFFF,
16'h021D, 16'hFFFF,
16'h021E, 16'hFFFF,
16'h021F, 16'hFFFF,
16'h0220, 16'hFFFF,
16'h0221, 16'hFFFF,
16'h0222, 16'hFFFF,
16'h0223, 16'hFFFF,
16'h0224, 16'hFFFF,
16'h0225, 16'hFFFF,
16'h0226, 16'hFFFF,
16'h0227, 16'hFFFF,
16'h0228, 16'hFFFF,
16'h0229, 16'hFFFF,
16'h022A, 16'hFFFF,
16'h022B, 16'hFFFF,
16'h022C, 16'hFFFF,
16'h022D, 16'hFFFF,
16'h022E, 16'hFFFF,
16'h022F, 16'hFFFF,
16'h0230, 16'hFFFF,
16'h0231, 16'hFFFF,
16'h0232, 16'hFFFF,
16'h0233, 16'hFFFF,
16'h0234, 16'hFFFF,
16'h0235, 16'hFFFF,
16'h0236, 16'hFFFF,
16'h0237, 16'hFFFF,
16'h0238, 16'hFFFF,
16'h0239, 16'hFFFF,
16'h023A, 16'hFFFF,
16'h023B, 16'hFFFF,
16'h023C, 16'hFFFF,
16'h023D, 16'hFFFF,
16'h023E, 16'hFFFF,
16'h023F, 16'hFFFF,
16'h0240, 16'hFFFF,
16'h0241, 16'hFFFF,
16'h0242, 16'hFFFF,
16'h0243, 16'hFFFF,
16'h0244, 16'hFFFF,
16'h0245, 16'hFFFF,
16'h0246, 16'hFFFF,
16'h0247, 16'hFFFF,
16'h0248, 16'hFFFF,
16'h0249, 16'hFFFF,
16'h024A, 16'hFFFF,
16'h024B, 16'hFFFF,
16'h024C, 16'hFFFF,
16'h024D, 16'hFFFF,
16'h024E, 16'hFFFF,
16'h024F, 16'hFFFF,
16'h0250, 16'hFFFF,
16'h0251, 16'hFFFF,
16'h0252, 16'hFFFF,
16'h0253, 16'hFFFF,
16'h0254, 16'hFFFF,
16'h0255, 16'hFFFF,
16'h0256, 16'hFFFF,
16'h0257, 16'hFFFF,
16'h0258, 16'hFFFF,
16'h0259, 16'hFFFF,
16'h025A, 16'hFFFF,
16'h025B, 16'hFFFF,
16'h025C, 16'hFFFF,
16'h025D, 16'hFFFF,
16'h025E, 16'hFFFF,
16'h025F, 16'hFFFF,
16'h0260, 16'hFFFF,
16'h0261, 16'hFFFF,
16'h0262, 16'hFFFF,
16'h0263, 16'hFFFF,
16'h0264, 16'hFFFF,
16'h0265, 16'hFFFF,
16'h0266, 16'hFFFF,
16'h0267, 16'hFFFF,
16'h0268, 16'hFFFF,
16'h0269, 16'hFFFF,
16'h026A, 16'hFFFF,
16'h026B, 16'hFFFF,
16'h026C, 16'hFFFF,
16'h026D, 16'hFFFF,
16'h026E, 16'hFFFF,
16'h026F, 16'hFFFF,
16'h0270, 16'hFFFF,
16'h0271, 16'hFFFF,
16'h0272, 16'hFFFF,
16'h0273, 16'hFFFF,
16'h0274, 16'hFFFF,
16'h0275, 16'hFFFF,
16'h0276, 16'hFFFF,
16'h0277, 16'hFFFF,
16'h0278, 16'hFFFF,
16'h0279, 16'hFFFF,
16'h027A, 16'hFFFF,
16'h027B, 16'hFFFF,
16'h027C, 16'hFFFF,
16'h027D, 16'hFFFF,
16'h027E, 16'hFFFF,
16'h027F, 16'hFFFF,
16'h0280, 16'hFFFF,
16'h0281, 16'hFFFF,
16'h0282, 16'hFFFF,
16'h0283, 16'hFFFF,
16'h0284, 16'hFFFF,
16'h0285, 16'hFFFF,
16'h0286, 16'hFFFF,
16'h0287, 16'hFFFF,
16'h0288, 16'hFFFF,
16'h0289, 16'hFFFF,
16'h028A, 16'hFFFF,
16'h028B, 16'hFFFF,
16'h028C, 16'hFFFF,
16'h028D, 16'hFFFF,
16'h028E, 16'hFFFF,
16'h028F, 16'hFFFF,
16'h0290, 16'hFFFF,
16'h0291, 16'hFFFF,
16'h0292, 16'hFFFF,
16'h0293, 16'hFFFF,
16'h0294, 16'hFFFF,
16'h0295, 16'hFFFF,
16'h0296, 16'hFFFF,
16'h0297, 16'hFFFF,
16'h0298, 16'hFFFF,
16'h0299, 16'hFFFF,
16'h029A, 16'hFFFF,
16'h029B, 16'hFFFF,
16'h029C, 16'hFFFF,
16'h029D, 16'hFFFF,
16'h029E, 16'hFFFF,
16'h029F, 16'hFFFF,
16'h02A0, 16'hFFFF,
16'h02A1, 16'hFFFF,
16'h02A2, 16'hFFFF,
16'h02A3, 16'hFFFF,
16'h02A4, 16'hFFFF,
16'h02A5, 16'hFFFF,
16'h02A6, 16'hFFFF,
16'h02A7, 16'hFFFF,
16'h02A8, 16'hFFFF,
16'h02A9, 16'hFFFF,
16'h02AA, 16'hFFFF,
16'h02AB, 16'hFFFF,
16'h02AC, 16'hFFFF,
16'h02AD, 16'hFFFF,
16'h02AE, 16'hFFFF,
16'h02AF, 16'hFFFF,
16'h02B0, 16'hFFFF,
16'h02B1, 16'hFFFF,
16'h02B2, 16'hFFFF,
16'h02B3, 16'hFFFF,
16'h02B4, 16'hFFFF,
16'h02B5, 16'hFFFF,
16'h02B6, 16'hFFFF,
16'h02B7, 16'hFFFF,
16'h02B8, 16'hFFFF,
16'h02B9, 16'hFFFF,
16'h02BA, 16'hFFFF,
16'h02BB, 16'hFFFF,
16'h02BC, 16'hFFFF,
16'h02BD, 16'hFFFF,
16'h02BE, 16'hFFFF,
16'h02BF, 16'hFFFF,
16'h02C0, 16'hFFFF,
16'h02C1, 16'hFFFF,
16'h02C2, 16'hFFFF,
16'h02C3, 16'hFFFF,
16'h02C4, 16'hFFFF,
16'h02C5, 16'hFFFF,
16'h02C6, 16'hFFFF,
16'h02C7, 16'hFFFF,
16'h02C8, 16'hFFFF,
16'h02C9, 16'hFFFF,
16'h02CA, 16'hFFFF,
16'h02CB, 16'hFFFF,
16'h02CC, 16'hFFFF,
16'h02CD, 16'hFFFF,
16'h02CE, 16'hFFFF,
16'h02CF, 16'hFFFF,
16'h02D0, 16'hFFFF,
16'h02D1, 16'hFFFF,
16'h02D2, 16'hFFFF,
16'h02D3, 16'hFFFF,
16'h02D4, 16'hFFFF,
16'h02D5, 16'hFFFF,
16'h02D6, 16'hFFFF,
16'h02D7, 16'hFFFF,
16'h02D8, 16'hFFFF,
16'h02D9, 16'hFFFF,
16'h02DA, 16'hFFFF,
16'h02DB, 16'hFFFF,
16'h02DC, 16'hFFFF,
16'h02DD, 16'hFFFF,
16'h02DE, 16'hFFFF,
16'h02DF, 16'hFFFF,
16'h02E0, 16'hFFFF,
16'h02E1, 16'hFFFF,
16'h02E2, 16'hFFFF,
16'h02E3, 16'hFFFF,
16'h02E4, 16'hFFFF,
16'h02E5, 16'hFFFF,
16'h02E6, 16'hFFFF,
16'h02E7, 16'hFFFF,
16'h02E8, 16'hFFFF,
16'h02E9, 16'hFFFF,
16'h02EA, 16'hFFFF,
16'h02EB, 16'hFFFF,
16'h02EC, 16'hFFFF,
16'h02ED, 16'hFFFF,
16'h02EE, 16'hFFFF,
16'h02EF, 16'hFFFF,
16'h02F0, 16'hFFFF,
16'h02F1, 16'hFFFF,
16'h02F2, 16'hFFFF,
16'h02F3, 16'hFFFF,
16'h02F4, 16'hFFFF,
16'h02F5, 16'hFFFF,
16'h02F6, 16'hFFFF,
16'h02F7, 16'hFFFF,
16'h02F8, 16'hFFFF,
16'h02F9, 16'hFFFF,
16'h02FA, 16'hFFFF,
16'h02FB, 16'hFFFF,
16'h02FC, 16'hFFFF,
16'h02FD, 16'hFFFF,
16'h02FE, 16'hFFFF,
16'h02FF, 16'hFFFF,
16'h0300, 16'hFFFF,
16'h0301, 16'hFFFF,
16'h0302, 16'hFFFF,
16'h0303, 16'hFFFF,
16'h0304, 16'hFFFF,
16'h0305, 16'hFFFF,
16'h0306, 16'hFFFF,
16'h0307, 16'hFFFF,
16'h0308, 16'hFFFF,
16'h0309, 16'hFFFF,
16'h030A, 16'hFFFF,
16'h030B, 16'hFFFF,
16'h030C, 16'hFFFF,
16'h030D, 16'hFFFF,
16'h030E, 16'hFFFF,
16'h030F, 16'hFFFF,
16'h0310, 16'hFFFF,
16'h0311, 16'hFFFF,
16'h0312, 16'hFFFF,
16'h0313, 16'hFFFF,
16'h0314, 16'hFFFF,
16'h0315, 16'hFFFF,
16'h0316, 16'hFFFF,
16'h0317, 16'hFFFF,
16'h0318, 16'hFFFF,
16'h0319, 16'hFFFF,
16'h031A, 16'hFFFF,
16'h031B, 16'hFFFF,
16'h031C, 16'hFFFF,
16'h031D, 16'hFFFF,
16'h031E, 16'hFFFF,
16'h031F, 16'hFFFF,
16'h0320, 16'hFFFF,
16'h0321, 16'hFFFF,
16'h0322, 16'hFFFF,
16'h0323, 16'hFFFF,
16'h0324, 16'hFFFF,
16'h0325, 16'hFFFF,
16'h0326, 16'hFFFF,
16'h0327, 16'hFFFF,
16'h0328, 16'hFFFF,
16'h0329, 16'hFFFF,
16'h032A, 16'hFFFF,
16'h032B, 16'hFFFF,
16'h032C, 16'hFFFF,
16'h032D, 16'hFFFF,
16'h032E, 16'hFFFF,
16'h032F, 16'hFFFF,
16'h0330, 16'hFFFF,
16'h0331, 16'hFFFF,
16'h0332, 16'hFFFF,
16'h0333, 16'hFFFF,
16'h0334, 16'hFFFF,
16'h0335, 16'hFFFF,
16'h0336, 16'hFFFF,
16'h0337, 16'hFFFF,
16'h0338, 16'hFFFF,
16'h0339, 16'hFFFF,
16'h033A, 16'hFFFF,
16'h033B, 16'hFFFF,
16'h033C, 16'hFFFF,
16'h033D, 16'hFFFF,
16'h033E, 16'hFFFF,
16'h033F, 16'hFFFF,
16'h0340, 16'hFFFF,
16'h0341, 16'hFFFF,
16'h0342, 16'hFFFF,
16'h0343, 16'hFFFF,
16'h0344, 16'hFFFF,
16'h0345, 16'hFFFF,
16'h0346, 16'hFFFF,
16'h0347, 16'hFFFF,
16'h0348, 16'hFFFF,
16'h0349, 16'hFFFF,
16'h034A, 16'hFFFF,
16'h034B, 16'hFFFF,
16'h034C, 16'hFFFF,
16'h034D, 16'hFFFF,
16'h034E, 16'hFFFF,
16'h034F, 16'hFFFF,
16'h0350, 16'hFFFF,
16'h0351, 16'hFFFF,
16'h0352, 16'hFFFF,
16'h0353, 16'hFFFF,
16'h0354, 16'hFFFF,
16'h0355, 16'hFFFF,
16'h0356, 16'hFFFF,
16'h0357, 16'hFFFF,
16'h0358, 16'hFFFF,
16'h0359, 16'hFFFF,
16'h035A, 16'hFFFF,
16'h035B, 16'hFFFF,
16'h035C, 16'hFFFF,
16'h035D, 16'hFFFF,
16'h035E, 16'hFFFF,
16'h035F, 16'hFFFF,
16'h0360, 16'hFFFF,
16'h0361, 16'hFFFF,
16'h0362, 16'hFFFF,
16'h0363, 16'hFFFF,
16'h0364, 16'hFFFF,
16'h0365, 16'hFFFF,
16'h0366, 16'hFFFF,
16'h0367, 16'hFFFF,
16'h0368, 16'hFFFF,
16'h0369, 16'hFFFF,
16'h036A, 16'hFFFF,
16'h036B, 16'hFFFF,
16'h036C, 16'hFFFF,
16'h036D, 16'hFFFF,
16'h036E, 16'hFFFF,
16'h036F, 16'hFFFF,
16'h0370, 16'hFFFF,
16'h0371, 16'hFFFF,
16'h0372, 16'hFFFF,
16'h0373, 16'hFFFF,
16'h0374, 16'hFFFF,
16'h0375, 16'hFFFF,
16'h0376, 16'hFFFF,
16'h0377, 16'hFFFF,
16'h0378, 16'hFFFF,
16'h0379, 16'hFFFF,
16'h037A, 16'hFFFF,
16'h037B, 16'hFFFF,
16'h037C, 16'hFFFF,
16'h037D, 16'hFFFF,
16'h037E, 16'hFFFF,
16'h037F, 16'hFFFF,
16'h0380, 16'hFFFF,
16'h0381, 16'hFFFF,
16'h0382, 16'hFFFF,
16'h0383, 16'hFFFF,
16'h0384, 16'hFFFF,
16'h0385, 16'hFFFF,
16'h0386, 16'hFFFF,
16'h0387, 16'hFFFF,
16'h0388, 16'hFFFF,
16'h0389, 16'hFFFF,
16'h038A, 16'hFFFF,
16'h038B, 16'hFFFF,
16'h038C, 16'hFFFF,
16'h038D, 16'hFFFF,
16'h038E, 16'hFFFF,
16'h038F, 16'hFFFF,
16'h0390, 16'hFFFF,
16'h0391, 16'hFFFF,
16'h0392, 16'hFFFF,
16'h0393, 16'hFFFF,
16'h0394, 16'hFFFF,
16'h0395, 16'hFFFF,
16'h0396, 16'hFFFF,
16'h0397, 16'hFFFF,
16'h0398, 16'hFFFF,
16'h0399, 16'hFFFF,
16'h039A, 16'hFFFF,
16'h039B, 16'hFFFF,
16'h039C, 16'hFFFF,
16'h039D, 16'hFFFF,
16'h039E, 16'hFFFF,
16'h039F, 16'hFFFF,
16'h03A0, 16'hFFFF,
16'h03A1, 16'hFFFF,
16'h03A2, 16'hFFFF,
16'h03A3, 16'hFFFF,
16'h03A4, 16'hFFFF,
16'h03A5, 16'hFFFF,
16'h03A6, 16'hFFFF,
16'h03A7, 16'hFFFF,
16'h03A8, 16'hFFFF,
16'h03A9, 16'hFFFF,
16'h03AA, 16'hFFFF,
16'h03AB, 16'hFFFF,
16'h03AC, 16'hFFFF,
16'h03AD, 16'hFFFF,
16'h03AE, 16'hFFFF,
16'h03AF, 16'hFFFF,
16'h03B0, 16'hFFFF,
16'h03B1, 16'hFFFF,
16'h03B2, 16'hFFFF,
16'h03B3, 16'hFFFF,
16'h03B4, 16'hFFFF,
16'h03B5, 16'hFFFF,
16'h03B6, 16'hFFFF,
16'h03B7, 16'hFFFF,
16'h03B8, 16'hFFFF,
16'h03B9, 16'hFFFF,
16'h03BA, 16'hFFFF,
16'h03BB, 16'hFFFF,
16'h03BC, 16'hFFFF,
16'h03BD, 16'hFFFF,
16'h03BE, 16'hFFFF,
16'h03BF, 16'hFFFF,
16'h03C0, 16'hFFFF,
16'h03C1, 16'hFFFF,
16'h03C2, 16'hFFFF,
16'h03C3, 16'hFFFF,
16'h03C4, 16'hFFFF,
16'h03C5, 16'hFFFF,
16'h03C6, 16'hFFFF,
16'h03C7, 16'hFFFF,
16'h03C8, 16'hFFFF,
16'h03C9, 16'hFFFF,
16'h03CA, 16'hFFFF,
16'h03CB, 16'hFFFF,
16'h03CC, 16'hFFFF,
16'h03CD, 16'hFFFF,
16'h03CE, 16'hFFFF,
16'h03CF, 16'hFFFF,
16'h03D0, 16'hFFFF,
16'h03D1, 16'hFFFF,
16'h03D2, 16'hFFFF,
16'h03D3, 16'hFFFF,
16'h03D4, 16'hFFFF,
16'h03D5, 16'hFFFF,
16'h03D6, 16'hFFFF,
16'h03D7, 16'hFFFF,
16'h03D8, 16'hFFFF,
16'h03D9, 16'hFFFF,
16'h03DA, 16'hFFFF,
16'h03DB, 16'hFFFF,
16'h03DC, 16'hFFFF,
16'h03DD, 16'hFFFF,
16'h03DE, 16'hFFFF,
16'h03DF, 16'hFFFF,
16'h03E0, 16'hFFFF,
16'h03E1, 16'hFFFF,
16'h03E2, 16'hFFFF,
16'h03E3, 16'hFFFF,
16'h03E4, 16'hFFFF,
16'h03E5, 16'hFFFF,
16'h03E6, 16'hFFFF,
16'h03E7, 16'hFFFF,
16'h03E8, 16'hFFFF,
16'h03E9, 16'hFFFF,
16'h03EA, 16'hFFFF,
16'h03EB, 16'hFFFF,
16'h03EC, 16'hFFFF,
16'h03ED, 16'hFFFF,
16'h03EE, 16'hFFFF,
16'h03EF, 16'hFFFF,
16'h03F0, 16'hFFFF,
16'h03F1, 16'hFFFF,
16'h03F2, 16'hFFFF,
16'h03F3, 16'hFFFF,
16'h03F4, 16'hFFFF,
16'h03F5, 16'hFFFF,
16'h03F6, 16'hFFFF,
16'h03F7, 16'hFFFF,
16'h03F8, 16'hFFFF,
16'h03F9, 16'hFFFF,
16'h03FA, 16'hFFFF,
16'h03FB, 16'hFFFF,
16'h03FC, 16'hFFFF,
16'h03FD, 16'hFFFF,
16'h03FE, 16'hFFFF,
16'h03FF, 16'hFFFF,
16'h0400, 16'hFFFF,
16'h0401, 16'hFFFF,
16'h0402, 16'hFFFF,
16'h0403, 16'hFFFF,
16'h0404, 16'hFFFF,
16'h0405, 16'hFFFF,
16'h0406, 16'hFFFF,
16'h0407, 16'hFFFF,
16'h0408, 16'hFFFF,
16'h0409, 16'hFFFF,
16'h040A, 16'hFFFF,
16'h040B, 16'hFFFF,
16'h040C, 16'hFFFF,
16'h040D, 16'hFFFF,
16'h040E, 16'hFFFF,
16'h040F, 16'hFFFF,
16'h0410, 16'hFFFF,
16'h0411, 16'hFFFF,
16'h0412, 16'hFFFF,
16'h0413, 16'hFFFF,
16'h0414, 16'hFFFF,
16'h0415, 16'hFFFF,
16'h0416, 16'hFFFF,
16'h0417, 16'hFFFF,
16'h0418, 16'hFFFF,
16'h0419, 16'hFFFF,
16'h041A, 16'hFFFF,
16'h041B, 16'hFFFF,
16'h041C, 16'hFFFF,
16'h041D, 16'hFFFF,
16'h041E, 16'hFFFF,
16'h041F, 16'hFFFF,
16'h0420, 16'hFFFF,
16'h0421, 16'hFFFF,
16'h0422, 16'hFFFF,
16'h0423, 16'hFFFF,
16'h0424, 16'hFFFF,
16'h0425, 16'hFFFF,
16'h0426, 16'hFFFF,
16'h0427, 16'hFFFF,
16'h0428, 16'hFFFF,
16'h0429, 16'hFFFF,
16'h042A, 16'hFFFF,
16'h042B, 16'hFFFF,
16'h042C, 16'hFFFF,
16'h042D, 16'hFFFF,
16'h042E, 16'hFFFF,
16'h042F, 16'hFFFF,
16'h0430, 16'hFFFF,
16'h0431, 16'hFFFF,
16'h0432, 16'hFFFF,
16'h0433, 16'hFFFF,
16'h0434, 16'hFFFF,
16'h0435, 16'hFFFF,
16'h0436, 16'hFFFF,
16'h0437, 16'hFFFF,
16'h0438, 16'hFFFF,
16'h0439, 16'hFFFF,
16'h043A, 16'hFFFF,
16'h043B, 16'hFFFF,
16'h043C, 16'hFFFF,
16'h043D, 16'hFFFF,
16'h043E, 16'hFFFF,
16'h043F, 16'hFFFF,
16'h0440, 16'hFFFF,
16'h0441, 16'hFFFF,
16'h0442, 16'hFFFF,
16'h0443, 16'hFFFF,
16'h0444, 16'hFFFF,
16'h0445, 16'hFFFF,
16'h0446, 16'hFFFF,
16'h0447, 16'hFFFF,
16'h0448, 16'hFFFF,
16'h0449, 16'hFFFF,
16'h044A, 16'hFFFF,
16'h044B, 16'hFFFF,
16'h044C, 16'hFFFF,
16'h044D, 16'hFFFF,
16'h044E, 16'hFFFF,
16'h044F, 16'hFFFF,
16'h0450, 16'hFFFF,
16'h0451, 16'hFFFF,
16'h0452, 16'hFFFF,
16'h0453, 16'hFFFF,
16'h0454, 16'hFFFF,
16'h0455, 16'hFFFF,
16'h0456, 16'hFFFF,
16'h0457, 16'hFFFF,
16'h0458, 16'hFFFF,
16'h0459, 16'hFFFF,
16'h045A, 16'hFFFF,
16'h045B, 16'hFFFF,
16'h045C, 16'hFFFF,
16'h045D, 16'hFFFF,
16'h045E, 16'hFFFF,
16'h045F, 16'hFFFF,
16'h0460, 16'hFFFF,
16'h0461, 16'hFFFF,
16'h0462, 16'hFFFF,
16'h0463, 16'hFFFF,
16'h0464, 16'hFFFF,
16'h0465, 16'hFFFF,
16'h0466, 16'hFFFF,
16'h0467, 16'hFFFF,
16'h0468, 16'hFFFF,
16'h0469, 16'hFFFF,
16'h046A, 16'hFFFF,
16'h046B, 16'hFFFF,
16'h046C, 16'hFFFF,
16'h046D, 16'hFFFF,
16'h046E, 16'hFFFF,
16'h046F, 16'hFFFF,
16'h0470, 16'hFFFF,
16'h0471, 16'hFFFF,
16'h0472, 16'hFFFF,
16'h0473, 16'hFFFF,
16'h0474, 16'hFFFF,
16'h0475, 16'hFFFF,
16'h0476, 16'hFFFF,
16'h0477, 16'hFFFF,
16'h0478, 16'hFFFF,
16'h0479, 16'hFFFF,
16'h047A, 16'hFFFF,
16'h047B, 16'hFFFF,
16'h047C, 16'hFFFF,
16'h047D, 16'hFFFF,
16'h047E, 16'hFFFF,
16'h047F, 16'hFFFF,
16'h0480, 16'hFFFF,
16'h0481, 16'hFFFF,
16'h0482, 16'hFFFF,
16'h0483, 16'hFFFF,
16'h0484, 16'hFFFF,
16'h0485, 16'hFFFF,
16'h0486, 16'hFFFF,
16'h0487, 16'hFFFF,
16'h0488, 16'hFFFF,
16'h0489, 16'hFFFF,
16'h048A, 16'hFFFF,
16'h048B, 16'hFFFF,
16'h048C, 16'hFFFF,
16'h048D, 16'hFFFF,
16'h048E, 16'hFFFF,
16'h048F, 16'hFFFF,
16'h0490, 16'hFFFF,
16'h0491, 16'hFFFF,
16'h0492, 16'hFFFF,
16'h0493, 16'hFFFF,
16'h0494, 16'hFFFF,
16'h0495, 16'hFFFF,
16'h0496, 16'hFFFF,
16'h0497, 16'hFFFF,
16'h0498, 16'hFFFF,
16'h0499, 16'hFFFF,
16'h049A, 16'hFFFF,
16'h049B, 16'hFFFF,
16'h049C, 16'hFFFF,
16'h049D, 16'hFFFF,
16'h049E, 16'hFFFF,
16'h049F, 16'hFFFF,
16'h04A0, 16'hFFFF,
16'h04A1, 16'hFFFF,
16'h04A2, 16'hFFFF,
16'h04A3, 16'hFFFF,
16'h04A4, 16'hFFFF,
16'h04A5, 16'hFFFF,
16'h04A6, 16'hFFFF,
16'h04A7, 16'hFFFF,
16'h04A8, 16'hFFFF,
16'h04A9, 16'hFFFF,
16'h04AA, 16'hFFFF,
16'h04AB, 16'hFFFF,
16'h04AC, 16'hFFFF,
16'h04AD, 16'hFFFF,
16'h04AE, 16'hFFFF,
16'h04AF, 16'hFFFF,
16'h04B0, 16'hFFFF,
16'h04B1, 16'hFFFF,
16'h04B2, 16'hFFFF,
16'h04B3, 16'hFFFF,
16'h04B4, 16'hFFFF,
16'h04B5, 16'hFFFF,
16'h04B6, 16'hFFFF,
16'h04B7, 16'hFFFF,
16'h04B8, 16'hFFFF,
16'h04B9, 16'hFFFF,
16'h04BA, 16'hFFFF,
16'h04BB, 16'hFFFF,
16'h04BC, 16'hFFFF,
16'h04BD, 16'hFFFF,
16'h04BE, 16'hFFFF,
16'h04BF, 16'hFFFF,
16'h04C0, 16'hFFFF,
16'h04C1, 16'hFFFF,
16'h04C2, 16'hFFFF,
16'h04C3, 16'hFFFF,
16'h04C4, 16'hFFFF,
16'h04C5, 16'hFFFF,
16'h04C6, 16'hFFFF,
16'h04C7, 16'hFFFF,
16'h04C8, 16'hFFFF,
16'h04C9, 16'hFFFF,
16'h04CA, 16'hFFFF,
16'h04CB, 16'hFFFF,
16'h04CC, 16'hFFFF,
16'h04CD, 16'hFFFF,
16'h04CE, 16'hFFFF,
16'h04CF, 16'hFFFF,
16'h04D0, 16'hFFFF,
16'h04D1, 16'hFFFF,
16'h04D2, 16'hFFFF,
16'h04D3, 16'hFFFF,
16'h04D4, 16'hFFFF,
16'h04D5, 16'hFFFF,
16'h04D6, 16'hFFFF,
16'h04D7, 16'hFFFF,
16'h04D8, 16'hFFFF,
16'h04D9, 16'hFFFF,
16'h04DA, 16'hFFFF,
16'h04DB, 16'hFFFF,
16'h04DC, 16'hFFFF,
16'h04DD, 16'hFFFF,
16'h04DE, 16'hFFFF,
16'h04DF, 16'hFFFF,
16'h04E0, 16'hFFFF,
16'h04E1, 16'hFFFF,
16'h04E2, 16'hFFFF,
16'h04E3, 16'hFFFF,
16'h04E4, 16'hFFFF,
16'h04E5, 16'hFFFF,
16'h04E6, 16'hFFFF,
16'h04E7, 16'hFFFF,
16'h04E8, 16'hFFFF,
16'h04E9, 16'hFFFF,
16'h04EA, 16'hFFFF,
16'h04EB, 16'hFFFF,
16'h04EC, 16'hFFFF,
16'h04ED, 16'hFFFF,
16'h04EE, 16'hFFFF,
16'h04EF, 16'hFFFF,
16'h04F0, 16'hFFFF,
16'h04F1, 16'hFFFF,
16'h04F2, 16'hFFFF,
16'h04F3, 16'hFFFF,
16'h04F4, 16'hFFFF,
16'h04F5, 16'hFFFF,
16'h04F6, 16'hFFFF,
16'h04F7, 16'hFFFF,
16'h04F8, 16'hFFFF,
16'h04F9, 16'hFFFF,
16'h04FA, 16'hFFFF,
16'h04FB, 16'hFFFF,
16'h04FC, 16'hFFFF,
16'h04FD, 16'hFFFF,
16'h04FE, 16'hFFFF,
16'h04FF, 16'hFFFF,
16'h0500, 16'hFFFF,
16'h0501, 16'hFFFF,
16'h0502, 16'hFFFF,
16'h0503, 16'hFFFF,
16'h0504, 16'hFFFF,
16'h0505, 16'hFFFF,
16'h0506, 16'hFFFF,
16'h0507, 16'hFFFF,
16'h0508, 16'hFFFF,
16'h0509, 16'hFFFF,
16'h050A, 16'hFFFF,
16'h050B, 16'hFFFF,
16'h050C, 16'hFFFF,
16'h050D, 16'hFFFF,
16'h050E, 16'hFFFF,
16'h050F, 16'hFFFF,
16'h0510, 16'hFFFF,
16'h0511, 16'hFFFF,
16'h0512, 16'hFFFF,
16'h0513, 16'hFFFF,
16'h0514, 16'hFFFF,
16'h0515, 16'hFFFF,
16'h0516, 16'hFFFF,
16'h0517, 16'hFFFF,
16'h0518, 16'hFFFF,
16'h0519, 16'hFFFF,
16'h051A, 16'hFFFF,
16'h051B, 16'hFFFF,
16'h051C, 16'hFFFF,
16'h051D, 16'hFFFF,
16'h051E, 16'hFFFF,
16'h051F, 16'hFFFF,
16'h0520, 16'hFFFF,
16'h0521, 16'hFFFF,
16'h0522, 16'hFFFF,
16'h0523, 16'hFFFF,
16'h0524, 16'hFFFF,
16'h0525, 16'hFFFF,
16'h0526, 16'hFFFF,
16'h0527, 16'hFFFF,
16'h0528, 16'hFFFF,
16'h0529, 16'hFFFF,
16'h052A, 16'hFFFF,
16'h052B, 16'hFFFF,
16'h052C, 16'hFFFF,
16'h052D, 16'hFFFF,
16'h052E, 16'hFFFF,
16'h052F, 16'hFFFF,
16'h0530, 16'hFFFF,
16'h0531, 16'hFFFF,
16'h0532, 16'hFFFF,
16'h0533, 16'hFFFF,
16'h0534, 16'hFFFF,
16'h0535, 16'hFFFF,
16'h0536, 16'hFFFF,
16'h0537, 16'hFFFF,
16'h0538, 16'hFFFF,
16'h0539, 16'hFFFF,
16'h053A, 16'hFFFF,
16'h053B, 16'hFFFF,
16'h053C, 16'hFFFF,
16'h053D, 16'hFFFF,
16'h053E, 16'hFFFF,
16'h053F, 16'hFFFF,
16'h0540, 16'hFFFF,
16'h0541, 16'hFFFF,
16'h0542, 16'hFFFF,
16'h0543, 16'hFFFF,
16'h0544, 16'hFFFF,
16'h0545, 16'hFFFF,
16'h0546, 16'hFFFF,
16'h0547, 16'hFFFF,
16'h0548, 16'hFFFF,
16'h0549, 16'hFFFF,
16'h054A, 16'hFFFF,
16'h054B, 16'hFFFF,
16'h054C, 16'hFFFF,
16'h054D, 16'hFFFF,
16'h054E, 16'hFFFF,
16'h054F, 16'hFFFF,
16'h0550, 16'hFFFF,
16'h0551, 16'hFFFF,
16'h0552, 16'hFFFF,
16'h0553, 16'hFFFF,
16'h0554, 16'hFFFF,
16'h0555, 16'hFFFF,
16'h0556, 16'hFFFF,
16'h0557, 16'hFFFF,
16'h0558, 16'hFFFF,
16'h0559, 16'hFFFF,
16'h055A, 16'hFFFF,
16'h055B, 16'hFFFF,
16'h055C, 16'hFFFF,
16'h055D, 16'hFFFF,
16'h055E, 16'hFFFF,
16'h055F, 16'hFFFF,
16'h0560, 16'hFFFF,
16'h0561, 16'hFFFF,
16'h0562, 16'hFFFF,
16'h0563, 16'hFFFF,
16'h0564, 16'hFFFF,
16'h0565, 16'hFFFF,
16'h0566, 16'hFFFF,
16'h0567, 16'hFFFF,
16'h0568, 16'hFFFF,
16'h0569, 16'hFFFF,
16'h056A, 16'hFFFF,
16'h056B, 16'hFFFF,
16'h056C, 16'hFFFF,
16'h056D, 16'hFFFF,
16'h056E, 16'hFFFF,
16'h056F, 16'hFFFF,
16'h0570, 16'hFFFF,
16'h0571, 16'hFFFF,
16'h0572, 16'hFFFF,
16'h0573, 16'hFFFF,
16'h0574, 16'hFFFF,
16'h0575, 16'hFFFF,
16'h0576, 16'hFFFF,
16'h0577, 16'hFFFF,
16'h0578, 16'hFFFF,
16'h0579, 16'hFFFF,
16'h057A, 16'hFFFF,
16'h057B, 16'hFFFF,
16'h057C, 16'hFFFF,
16'h057D, 16'hFFFF,
16'h057E, 16'hFFFF,
16'h057F, 16'hFFFF,
16'h0580, 16'hFFFF,
16'h0581, 16'hFFFF,
16'h0582, 16'hFFFF,
16'h0583, 16'hFFFF,
16'h0584, 16'hFFFF,
16'h0585, 16'hFFFF,
16'h0586, 16'hFFFF,
16'h0587, 16'hFFFF,
16'h0588, 16'hFFFF,
16'h0589, 16'hFFFF,
16'h058A, 16'hFFFF,
16'h058B, 16'hFFFF,
16'h058C, 16'hFFFF,
16'h058D, 16'hFFFF,
16'h058E, 16'hFFFF,
16'h058F, 16'hFFFF,
16'h0590, 16'hFFFF,
16'h0591, 16'hFFFF,
16'h0592, 16'hFFFF,
16'h0593, 16'hFFFF,
16'h0594, 16'hFFFF,
16'h0595, 16'hFFFF,
16'h0596, 16'hFFFF,
16'h0597, 16'hFFFF,
16'h0598, 16'hFFFF,
16'h0599, 16'hFFFF,
16'h059A, 16'hFFFF,
16'h059B, 16'hFFFF,
16'h059C, 16'hFFFF,
16'h059D, 16'hFFFF,
16'h059E, 16'hFFFF,
16'h059F, 16'hFFFF,
16'h05A0, 16'hFFFF,
16'h05A1, 16'hFFFF,
16'h05A2, 16'hFFFF,
16'h05A3, 16'hFFFF,
16'h05A4, 16'hFFFF,
16'h05A5, 16'hFFFF,
16'h05A6, 16'hFFFF,
16'h05A7, 16'hFFFF,
16'h05A8, 16'hFFFF,
16'h05A9, 16'hFFFF,
16'h05AA, 16'hFFFF,
16'h05AB, 16'hFFFF,
16'h05AC, 16'hFFFF,
16'h05AD, 16'hFFFF,
16'h05AE, 16'hFFFF,
16'h05AF, 16'hFFFF,
16'h05B0, 16'hFFFF,
16'h05B1, 16'hFFFF,
16'h05B2, 16'hFFFF,
16'h05B3, 16'hFFFF,
16'h05B4, 16'hFFFF,
16'h05B5, 16'hFFFF,
16'h05B6, 16'hFFFF,
16'h05B7, 16'hFFFF,
16'h05B8, 16'hFFFF,
16'h05B9, 16'hFFFF,
16'h05BA, 16'hFFFF,
16'h05BB, 16'hFFFF,
16'h05BC, 16'hFFFF,
16'h05BD, 16'hFFFF,
16'h05BE, 16'hFFFF,
16'h05BF, 16'hFFFF,
16'h05C0, 16'hFFFF,
16'h05C1, 16'hFFFF,
16'h05C2, 16'hFFFF,
16'h05C3, 16'hFFFF,
16'h05C4, 16'hFFFF,
16'h05C5, 16'hFFFF,
16'h05C6, 16'hFFFF,
16'h05C7, 16'hFFFF,
16'h05C8, 16'hFFFF,
16'h05C9, 16'hFFFF,
16'h05CA, 16'hFFFF,
16'h05CB, 16'hFFFF,
16'h05CC, 16'hFFFF,
16'h05CD, 16'hFFFF,
16'h05CE, 16'hFFFF,
16'h05CF, 16'hFFFF,
16'h05D0, 16'hFFFF,
16'h05D1, 16'hFFFF,
16'h05D2, 16'hFFFF,
16'h05D3, 16'hFFFF,
16'h05D4, 16'hFFFF,
16'h05D5, 16'hFFFF,
16'h05D6, 16'hFFFF,
16'h05D7, 16'hFFFF,
16'h05D8, 16'hFFFF,
16'h05D9, 16'hFFFF,
16'h05DA, 16'hFFFF,
16'h05DB, 16'hFFFF,
16'h05DC, 16'hFFFF,
16'h05DD, 16'hFFFF,
16'h05DE, 16'hFFFF,
16'h05DF, 16'hFFFF,
16'h05E0, 16'hFFFF,
16'h05E1, 16'hFFFF,
16'h05E2, 16'hFFFF,
16'h05E3, 16'hFFFF,
16'h05E4, 16'hFFFF,
16'h05E5, 16'hFFFF,
16'h05E6, 16'hFFFF,
16'h05E7, 16'hFFFF,
16'h05E8, 16'hFFFF,
16'h05E9, 16'hFFFF,
16'h05EA, 16'hFFFF,
16'h05EB, 16'hFFFF,
16'h05EC, 16'hFFFF,
16'h05ED, 16'hFFFF,
16'h05EE, 16'hFFFF,
16'h05EF, 16'hFFFF,
16'h05F0, 16'hFFFF,
16'h05F1, 16'hFFFF,
16'h05F2, 16'hFFFF,
16'h05F3, 16'hFFFF,
16'h05F4, 16'hFFFF,
16'h05F5, 16'hFFFF,
16'h05F6, 16'hFFFF,
16'h05F7, 16'hFFFF,
16'h05F8, 16'hFFFF,
16'h05F9, 16'hFFFF,
16'h05FA, 16'hFFFF,
16'h05FB, 16'hFFFF,
16'h05FC, 16'hFFFF,
16'h05FD, 16'hFFFF,
16'h05FE, 16'hFFFF,
16'h05FF, 16'hFFFF,
16'h0600, 16'hFFFF,
16'h0601, 16'hFFFF,
16'h0602, 16'hFFFF,
16'h0603, 16'hFFFF,
16'h0604, 16'hFFFF,
16'h0605, 16'hFFFF,
16'h0606, 16'hFFFF,
16'h0607, 16'hFFFF,
16'h0608, 16'hFFFF,
16'h0609, 16'hFFFF,
16'h060A, 16'hFFFF,
16'h060B, 16'hFFFF,
16'h060C, 16'hFFFF,
16'h060D, 16'hFFFF,
16'h060E, 16'hFFFF,
16'h060F, 16'hFFFF,
16'h0610, 16'hFFFF,
16'h0611, 16'hFFFF,
16'h0612, 16'hFFFF,
16'h0613, 16'hFFFF,
16'h0614, 16'hFFFF,
16'h0615, 16'hFFFF,
16'h0616, 16'hFFFF,
16'h0617, 16'hFFFF,
16'h0618, 16'hFFFF,
16'h0619, 16'hFFFF,
16'h061A, 16'hFFFF,
16'h061B, 16'hFFFF,
16'h061C, 16'hFFFF,
16'h061D, 16'hFFFF,
16'h061E, 16'hFFFF,
16'h061F, 16'hFFFF,
16'h0620, 16'hFFFF,
16'h0621, 16'hFFFF,
16'h0622, 16'hFFFF,
16'h0623, 16'hFFFF,
16'h0624, 16'hFFFF,
16'h0625, 16'hFFFF,
16'h0626, 16'hFFFF,
16'h0627, 16'hFFFF,
16'h0628, 16'hFFFF,
16'h0629, 16'hFFFF,
16'h062A, 16'hFFFF,
16'h062B, 16'hFFFF,
16'h062C, 16'hFFFF,
16'h062D, 16'hFFFF,
16'h062E, 16'hFFFF,
16'h062F, 16'hFFFF,
16'h0630, 16'hFFFF,
16'h0631, 16'hFFFF,
16'h0632, 16'hFFFF,
16'h0633, 16'hFFFF,
16'h0634, 16'hFFFF,
16'h0635, 16'hFFFF,
16'h0636, 16'hFFFF,
16'h0637, 16'hFFFF,
16'h0638, 16'hFFFF,
16'h0639, 16'hFFFF,
16'h063A, 16'hFFFF,
16'h063B, 16'hFFFF,
16'h063C, 16'hFFFF,
16'h063D, 16'hFFFF,
16'h063E, 16'hFFFF,
16'h063F, 16'hFFFF,
16'h0640, 16'hFFFF,
16'h0641, 16'hFFFF,
16'h0642, 16'hFFFF,
16'h0643, 16'hFFFF,
16'h0644, 16'hFFFF,
16'h0645, 16'hFFFF,
16'h0646, 16'hFFFF,
16'h0647, 16'hFFFF,
16'h0648, 16'hFFFF,
16'h0649, 16'hFFFF,
16'h064A, 16'hFFFF,
16'h064B, 16'hFFFF,
16'h064C, 16'hFFFF,
16'h064D, 16'hFFFF,
16'h064E, 16'hFFFF,
16'h064F, 16'hFFFF,
16'h0650, 16'hFFFF,
16'h0651, 16'hFFFF,
16'h0652, 16'hFFFF,
16'h0653, 16'hFFFF,
16'h0654, 16'hFFFF,
16'h0655, 16'hFFFF,
16'h0656, 16'hFFFF,
16'h0657, 16'hFFFF,
16'h0658, 16'hFFFF,
16'h0659, 16'hFFFF,
16'h065A, 16'hFFFF,
16'h065B, 16'hFFFF,
16'h065C, 16'hFFFF,
16'h065D, 16'hFFFF,
16'h065E, 16'hFFFF,
16'h065F, 16'hFFFF,
16'h0660, 16'hFFFF,
16'h0661, 16'hFFFF,
16'h0662, 16'hFFFF,
16'h0663, 16'hFFFF,
16'h0664, 16'hFFFF,
16'h0665, 16'hFFFF,
16'h0666, 16'hFFFF,
16'h0667, 16'hFFFF,
16'h0668, 16'hFFFF,
16'h0669, 16'hFFFF,
16'h066A, 16'hFFFF,
16'h066B, 16'hFFFF,
16'h066C, 16'hFFFF,
16'h066D, 16'hFFFF,
16'h066E, 16'hFFFF,
16'h066F, 16'hFFFF,
16'h0670, 16'hFFFF,
16'h0671, 16'hFFFF,
16'h0672, 16'hFFFF,
16'h0673, 16'hFFFF,
16'h0674, 16'hFFFF,
16'h0675, 16'hFFFF,
16'h0676, 16'hFFFF,
16'h0677, 16'hFFFF,
16'h0678, 16'hFFFF,
16'h0679, 16'hFFFF,
16'h067A, 16'hFFFF,
16'h067B, 16'hFFFF,
16'h067C, 16'hFFFF,
16'h067D, 16'hFFFF,
16'h067E, 16'hFFFF,
16'h067F, 16'hFFFF,
16'h0680, 16'hFFFF,
16'h0681, 16'hFFFF,
16'h0682, 16'hFFFF,
16'h0683, 16'hFFFF,
16'h0684, 16'hFFFF,
16'h0685, 16'hFFFF,
16'h0686, 16'hFFFF,
16'h0687, 16'hFFFF,
16'h0688, 16'hFFFF,
16'h0689, 16'hFFFF,
16'h068A, 16'hFFFF,
16'h068B, 16'hFFFF,
16'h068C, 16'hFFFF,
16'h068D, 16'hFFFF,
16'h068E, 16'hFFFF,
16'h068F, 16'hFFFF,
16'h0690, 16'hFFFF,
16'h0691, 16'hFFFF,
16'h0692, 16'hFFFF,
16'h0693, 16'hFFFF,
16'h0694, 16'hFFFF,
16'h0695, 16'hFFFF,
16'h0696, 16'hFFFF,
16'h0697, 16'hFFFF,
16'h0698, 16'hFFFF,
16'h0699, 16'hFFFF,
16'h069A, 16'hFFFF,
16'h069B, 16'hFFFF,
16'h069C, 16'hFFFF,
16'h069D, 16'hFFFF,
16'h069E, 16'hFFFF,
16'h069F, 16'hFFFF,
16'h06A0, 16'hFFFF,
16'h06A1, 16'hFFFF,
16'h06A2, 16'hFFFF,
16'h06A3, 16'hFFFF,
16'h06A4, 16'hFFFF,
16'h06A5, 16'hFFFF,
16'h06A6, 16'hFFFF,
16'h06A7, 16'hFFFF,
16'h06A8, 16'hFFFF,
16'h06A9, 16'hFFFF,
16'h06AA, 16'hFFFF,
16'h06AB, 16'hFFFF,
16'h06AC, 16'hFFFF,
16'h06AD, 16'hFFFF,
16'h06AE, 16'hFFFF,
16'h06AF, 16'hFFFF,
16'h06B0, 16'hFFFF,
16'h06B1, 16'hFFFF,
16'h06B2, 16'hFFFF,
16'h06B3, 16'hFFFF,
16'h06B4, 16'hFFFF,
16'h06B5, 16'hFFFF,
16'h06B6, 16'hFFFF,
16'h06B7, 16'hFFFF,
16'h06B8, 16'hFFFF,
16'h06B9, 16'hFFFF,
16'h06BA, 16'hFFFF,
16'h06BB, 16'hFFFF,
16'h06BC, 16'hFFFF,
16'h06BD, 16'hFFFF,
16'h06BE, 16'hFFFF,
16'h06BF, 16'hFFFF,
16'h06C0, 16'hFFFF,
16'h06C1, 16'hFFFF,
16'h06C2, 16'hFFFF,
16'h06C3, 16'hFFFF,
16'h06C4, 16'hFFFF,
16'h06C5, 16'hFFFF,
16'h06C6, 16'hFFFF,
16'h06C7, 16'hFFFF,
16'h06C8, 16'hFFFF,
16'h06C9, 16'hFFFF,
16'h06CA, 16'hFFFF,
16'h06CB, 16'hFFFF,
16'h06CC, 16'hFFFF,
16'h06CD, 16'hFFFF,
16'h06CE, 16'hFFFF,
16'h06CF, 16'hFFFF,
16'h06D0, 16'hFFFF,
16'h06D1, 16'hFFFF,
16'h06D2, 16'hFFFF,
16'h06D3, 16'hFFFF,
16'h06D4, 16'hFFFF,
16'h06D5, 16'hFFFF,
16'h06D6, 16'hFFFF,
16'h06D7, 16'hFFFF,
16'h06D8, 16'hFFFF,
16'h06D9, 16'hFFFF,
16'h06DA, 16'hFFFF,
16'h06DB, 16'hFFFF,
16'h06DC, 16'hFFFF,
16'h06DD, 16'hFFFF,
16'h06DE, 16'hFFFF,
16'h06DF, 16'hFFFF,
16'h06E0, 16'hFFFF,
16'h06E1, 16'hFFFF,
16'h06E2, 16'hFFFF,
16'h06E3, 16'hFFFF,
16'h06E4, 16'hFFFF,
16'h06E5, 16'hFFFF,
16'h06E6, 16'hFFFF,
16'h06E7, 16'hFFFF,
16'h06E8, 16'hFFFF,
16'h06E9, 16'hFFFF,
16'h06EA, 16'hFFFF,
16'h06EB, 16'hFFFF,
16'h06EC, 16'hFFFF,
16'h06ED, 16'hFFFF,
16'h06EE, 16'hFFFF,
16'h06EF, 16'hFFFF,
16'h06F0, 16'hFFFF,
16'h06F1, 16'hFFFF,
16'h06F2, 16'hFFFF,
16'h06F3, 16'hFFFF,
16'h06F4, 16'hFFFF,
16'h06F5, 16'hFFFF,
16'h06F6, 16'hFFFF,
16'h06F7, 16'hFFFF,
16'h06F8, 16'hFFFF,
16'h06F9, 16'hFFFF,
16'h06FA, 16'hFFFF,
16'h06FB, 16'hFFFF,
16'h06FC, 16'hFFFF,
16'h06FD, 16'hFFFF,
16'h06FE, 16'hFFFF,
16'h06FF, 16'hFFFF,
16'h0700, 16'hFFFF,
16'h0701, 16'hFFFF,
16'h0702, 16'hFFFF,
16'h0703, 16'hFFFF,
16'h0704, 16'hFFFF,
16'h0705, 16'hFFFF,
16'h0706, 16'hFFFF,
16'h0707, 16'hFFFF,
16'h0708, 16'hFFFF,
16'h0709, 16'hFFFF,
16'h070A, 16'hFFFF,
16'h070B, 16'hFFFF,
16'h070C, 16'hFFFF,
16'h070D, 16'hFFFF,
16'h070E, 16'hFFFF,
16'h070F, 16'hFFFF,
16'h0710, 16'hFFFF,
16'h0711, 16'hFFFF,
16'h0712, 16'hFFFF,
16'h0713, 16'hFFFF,
16'h0714, 16'hFFFF,
16'h0715, 16'hFFFF,
16'h0716, 16'hFFFF,
16'h0717, 16'hFFFF,
16'h0718, 16'hFFFF,
16'h0719, 16'hFFFF,
16'h071A, 16'hFFFF,
16'h071B, 16'hFFFF,
16'h071C, 16'hFFFF,
16'h071D, 16'hFFFF,
16'h071E, 16'hFFFF,
16'h071F, 16'hFFFF,
16'h0720, 16'hFFFF,
16'h0721, 16'hFFFF,
16'h0722, 16'hFFFF,
16'h0723, 16'hFFFF,
16'h0724, 16'hFFFF,
16'h0725, 16'hFFFF,
16'h0726, 16'hFFFF,
16'h0727, 16'hFFFF,
16'h0728, 16'hFFFF,
16'h0729, 16'hFFFF,
16'h072A, 16'hFFFF,
16'h072B, 16'hFFFF,
16'h072C, 16'hFFFF,
16'h072D, 16'hFFFF,
16'h072E, 16'hFFFF,
16'h072F, 16'hFFFF,
16'h0730, 16'hFFFF,
16'h0731, 16'hFFFF,
16'h0732, 16'hFFFF,
16'h0733, 16'hFFFF,
16'h0734, 16'hFFFF,
16'h0735, 16'hFFFF,
16'h0736, 16'hFFFF,
16'h0737, 16'hFFFF,
16'h0738, 16'hFFFF,
16'h0739, 16'hFFFF,
16'h073A, 16'hFFFF,
16'h073B, 16'hFFFF,
16'h073C, 16'hFFFF,
16'h073D, 16'hFFFF,
16'h073E, 16'hFFFF,
16'h073F, 16'hFFFF,
16'h0740, 16'hFFFF,
16'h0741, 16'hFFFF,
16'h0742, 16'hFFFF,
16'h0743, 16'hFFFF,
16'h0744, 16'hFFFF,
16'h0745, 16'hFFFF,
16'h0746, 16'hFFFF,
16'h0747, 16'hFFFF,
16'h0748, 16'hFFFF,
16'h0749, 16'hFFFF,
16'h074A, 16'hFFFF,
16'h074B, 16'hFFFF,
16'h074C, 16'hFFFF,
16'h074D, 16'hFFFF,
16'h074E, 16'hFFFF,
16'h074F, 16'hFFFF,
16'h0750, 16'hFFFF,
16'h0751, 16'hFFFF,
16'h0752, 16'hFFFF,
16'h0753, 16'hFFFF,
16'h0754, 16'hFFFF,
16'h0755, 16'hFFFF,
16'h0756, 16'hFFFF,
16'h0757, 16'hFFFF,
16'h0758, 16'hFFFF,
16'h0759, 16'hFFFF,
16'h075A, 16'hFFFF,
16'h075B, 16'hFFFF,
16'h075C, 16'hFFFF,
16'h075D, 16'hFFFF,
16'h075E, 16'hFFFF,
16'h075F, 16'hFFFF,
16'h0760, 16'hFFFF,
16'h0761, 16'hFFFF,
16'h0762, 16'hFFFF,
16'h0763, 16'hFFFF,
16'h0764, 16'hFFFF,
16'h0765, 16'hFFFF,
16'h0766, 16'hFFFF,
16'h0767, 16'hFFFF,
16'h0768, 16'hFFFF,
16'h0769, 16'hFFFF,
16'h076A, 16'hFFFF,
16'h076B, 16'hFFFF,
16'h076C, 16'hFFFF,
16'h076D, 16'hFFFF,
16'h076E, 16'hFFFF,
16'h076F, 16'hFFFF,
16'h0770, 16'hFFFF,
16'h0771, 16'hFFFF,
16'h0772, 16'hFFFF,
16'h0773, 16'hFFFF,
16'h0774, 16'hFFFF,
16'h0775, 16'hFFFF,
16'h0776, 16'hFFFF,
16'h0777, 16'hFFFF,
16'h0778, 16'hFFFF,
16'h0779, 16'hFFFF,
16'h077A, 16'hFFFF,
16'h077B, 16'hFFFF,
16'h077C, 16'hFFFF,
16'h077D, 16'hFFFF,
16'h077E, 16'hFFFF,
16'h077F, 16'hFFFF,
16'h0780, 16'hFFFF,
16'h0781, 16'hFFFF,
16'h0782, 16'hFFFF,
16'h0783, 16'hFFFF,
16'h0784, 16'hFFFF,
16'h0785, 16'hFFFF,
16'h0786, 16'hFFFF,
16'h0787, 16'hFFFF,
16'h0788, 16'hFFFF,
16'h0789, 16'hFFFF,
16'h078A, 16'hFFFF,
16'h078B, 16'hFFFF,
16'h078C, 16'hFFFF,
16'h078D, 16'hFFFF,
16'h078E, 16'hFFFF,
16'h078F, 16'hFFFF,
16'h0790, 16'hFFFF,
16'h0791, 16'hFFFF,
16'h0792, 16'hFFFF,
16'h0793, 16'hFFFF,
16'h0794, 16'hFFFF,
16'h0795, 16'hFFFF,
16'h0796, 16'hFFFF,
16'h0797, 16'hFFFF,
16'h0798, 16'hFFFF,
16'h0799, 16'hFFFF,
16'h079A, 16'hFFFF,
16'h079B, 16'hFFFF,
16'h079C, 16'hFFFF,
16'h079D, 16'hFFFF,
16'h079E, 16'hFFFF,
16'h079F, 16'hFFFF,
16'h07A0, 16'hFFFF,
16'h07A1, 16'hFFFF,
16'h07A2, 16'hFFFF,
16'h07A3, 16'hFFFF,
16'h07A4, 16'hFFFF,
16'h07A5, 16'hFFFF,
16'h07A6, 16'hFFFF,
16'h07A7, 16'hFFFF,
16'h07A8, 16'hFFFF,
16'h07A9, 16'hFFFF,
16'h07AA, 16'hFFFF,
16'h07AB, 16'hFFFF,
16'h07AC, 16'hFFFF,
16'h07AD, 16'hFFFF,
16'h07AE, 16'hFFFF,
16'h07AF, 16'hFFFF,
16'h07B0, 16'hFFFF,
16'h07B1, 16'hFFFF,
16'h07B2, 16'hFFFF,
16'h07B3, 16'hFFFF,
16'h07B4, 16'hFFFF,
16'h07B5, 16'hFFFF,
16'h07B6, 16'hFFFF,
16'h07B7, 16'hFFFF,
16'h07B8, 16'hFFFF,
16'h07B9, 16'hFFFF,
16'h07BA, 16'hFFFF,
16'h07BB, 16'hFFFF,
16'h07BC, 16'hFFFF,
16'h07BD, 16'hFFFF,
16'h07BE, 16'hFFFF,
16'h07BF, 16'hFFFF,
16'h07C0, 16'hFFFF,
16'h07C1, 16'hFFFF,
16'h07C2, 16'hFFFF,
16'h07C3, 16'hFFFF,
16'h07C4, 16'hFFFF,
16'h07C5, 16'hFFFF,
16'h07C6, 16'hFFFF,
16'h07C7, 16'hFFFF,
16'h07C8, 16'hFFFF,
16'h07C9, 16'hFFFF,
16'h07CA, 16'hFFFF,
16'h07CB, 16'hFFFF,
16'h07CC, 16'hFFFF,
16'h07CD, 16'hFFFF,
16'h07CE, 16'hFFFF,
16'h07CF, 16'hFFFF,
16'h07D0, 16'hFFFF,
16'h07D1, 16'hFFFF,
16'h07D2, 16'hFFFF,
16'h07D3, 16'hFFFF,
16'h07D4, 16'hFFFF,
16'h07D5, 16'hFFFF,
16'h07D6, 16'hFFFF,
16'h07D7, 16'hFFFF,
16'h07D8, 16'hFFFF,
16'h07D9, 16'hFFFF,
16'h07DA, 16'hFFFF,
16'h07DB, 16'hFFFF,
16'h07DC, 16'hFFFF,
16'h07DD, 16'hFFFF,
16'h07DE, 16'hFFFF,
16'h07DF, 16'hFFFF,
16'h07E0, 16'hFFFF,
16'h07E1, 16'hFFFF,
16'h07E2, 16'hFFFF,
16'h07E3, 16'hFFFF,
16'h07E4, 16'hFFFF,
16'h07E5, 16'hFFFF,
16'h07E6, 16'hFFFF,
16'h07E7, 16'hFFFF,
16'h07E8, 16'hFFFF,
16'h07E9, 16'hFFFF,
16'h07EA, 16'hFFFF,
16'h07EB, 16'hFFFF,
16'h07EC, 16'hFFFF,
16'h07ED, 16'hFFFF,
16'h07EE, 16'hFFFF,
16'h07EF, 16'hFFFF,
16'h07F0, 16'hFFFF,
16'h07F1, 16'hFFFF,
16'h07F2, 16'hFFFF,
16'h07F3, 16'hFFFF,
16'h07F4, 16'hFFFF,
16'h07F5, 16'hFFFF,
16'h07F6, 16'hFFFF,
16'h07F7, 16'hFFFF,
16'h07F8, 16'hFFFF,
16'h07F9, 16'hFFFF,
16'h07FA, 16'hFFFF,
16'h07FB, 16'hFFFF,
16'h07FC, 16'hFFFF,
16'h07FD, 16'hFFFF,
16'h07FE, 16'hFFFF,
16'h07FF, 16'hFFFF,
16'h0800, 16'hFFFF,
16'h0801, 16'hFFFF,
16'h0802, 16'hFFFF,
16'h0803, 16'hFFFF,
16'h0804, 16'hFFFF,
16'h0805, 16'hFFFF,
16'h0806, 16'hFFFF,
16'h0807, 16'hFFFF,
16'h0808, 16'hFFFF,
16'h0809, 16'hFFFF,
16'h080A, 16'hFFFF,
16'h080B, 16'hFFFF,
16'h080C, 16'hFFFF,
16'h080D, 16'hFFFF,
16'h080E, 16'hFFFF,
16'h080F, 16'hFFFF,
16'h0810, 16'hFFFF,
16'h0811, 16'hFFFF,
16'h0812, 16'hFFFF,
16'h0813, 16'hFFFF,
16'h0814, 16'hFFFF,
16'h0815, 16'hFFFF,
16'h0816, 16'hFFFF,
16'h0817, 16'hFFFF,
16'h0818, 16'hFFFF,
16'h0819, 16'hFFFF,
16'h081A, 16'hFFFF,
16'h081B, 16'hFFFF,
16'h081C, 16'hFFFF,
16'h081D, 16'hFFFF,
16'h081E, 16'hFFFF,
16'h081F, 16'hFFFF,
16'h0820, 16'hFFFF,
16'h0821, 16'hFFFF,
16'h0822, 16'hFFFF,
16'h0823, 16'hFFFF,
16'h0824, 16'hFFFF,
16'h0825, 16'hFFFF,
16'h0826, 16'hFFFF,
16'h0827, 16'hFFFF,
16'h0828, 16'hFFFF,
16'h0829, 16'hFFFF,
16'h082A, 16'hFFFF,
16'h082B, 16'hFFFF,
16'h082C, 16'hFFFF,
16'h082D, 16'hFFFF,
16'h082E, 16'hFFFF,
16'h082F, 16'hFFFF,
16'h0830, 16'hFFFF,
16'h0831, 16'hFFFF,
16'h0832, 16'hFFFF,
16'h0833, 16'hFFFF,
16'h0834, 16'hFFFF,
16'h0835, 16'hFFFF,
16'h0836, 16'hFFFF,
16'h0837, 16'hFFFF,
16'h0838, 16'hFFFF,
16'h0839, 16'hFFFF,
16'h083A, 16'hFFFF,
16'h083B, 16'hFFFF,
16'h083C, 16'hFFFF,
16'h083D, 16'hFFFF,
16'h083E, 16'hFFFF,
16'h083F, 16'hFFFF,
16'h0840, 16'hFFFF,
16'h0841, 16'hFFFF,
16'h0842, 16'hFFFF,
16'h0843, 16'hFFFF,
16'h0844, 16'hFFFF,
16'h0845, 16'hFFFF,
16'h0846, 16'hFFFF,
16'h0847, 16'hFFFF,
16'h0848, 16'hFFFF,
16'h0849, 16'hFFFF,
16'h084A, 16'hFFFF,
16'h084B, 16'hFFFF,
16'h084C, 16'hFFFF,
16'h084D, 16'hFFFF,
16'h084E, 16'hFFFF,
16'h084F, 16'hFFFF,
16'h0850, 16'hFFFF,
16'h0851, 16'hFFFF,
16'h0852, 16'hFFFF,
16'h0853, 16'hFFFF,
16'h0854, 16'hFFFF,
16'h0855, 16'hFFFF,
16'h0856, 16'hFFFF,
16'h0857, 16'hFFFF,
16'h0858, 16'hFFFF,
16'h0859, 16'hFFFF,
16'h085A, 16'hFFFF,
16'h085B, 16'hFFFF,
16'h085C, 16'hFFFF,
16'h085D, 16'hFFFF,
16'h085E, 16'hFFFF,
16'h085F, 16'hFFFF,
16'h0860, 16'hFFFF,
16'h0861, 16'hFFFF,
16'h0862, 16'hFFFF,
16'h0863, 16'hFFFF,
16'h0864, 16'hFFFF,
16'h0865, 16'hFFFF,
16'h0866, 16'hFFFF,
16'h0867, 16'hFFFF,
16'h0868, 16'hFFFF,
16'h0869, 16'hFFFF,
16'h086A, 16'hFFFF,
16'h086B, 16'hFFFF,
16'h086C, 16'hFFFF,
16'h086D, 16'hFFFF,
16'h086E, 16'hFFFF,
16'h086F, 16'hFFFF,
16'h0870, 16'hFFFF,
16'h0871, 16'hFFFF,
16'h0872, 16'hFFFF,
16'h0873, 16'hFFFF,
16'h0874, 16'hFFFF,
16'h0875, 16'hFFFF,
16'h0876, 16'hFFFF,
16'h0877, 16'hFFFF,
16'h0878, 16'hFFFF,
16'h0879, 16'hFFFF,
16'h087A, 16'hFFFF,
16'h087B, 16'hFFFF,
16'h087C, 16'hFFFF,
16'h087D, 16'hFFFF,
16'h087E, 16'hFFFF,
16'h087F, 16'hFFFF,
16'h0880, 16'hFFFF,
16'h0881, 16'hFFFF,
16'h0882, 16'hFFFF,
16'h0883, 16'hFFFF,
16'h0884, 16'hFFFF,
16'h0885, 16'hFFFF,
16'h0886, 16'hFFFF,
16'h0887, 16'hFFFF,
16'h0888, 16'hFFFF,
16'h0889, 16'hFFFF,
16'h088A, 16'hFFFF,
16'h088B, 16'hFFFF,
16'h088C, 16'hFFFF,
16'h088D, 16'hFFFF,
16'h088E, 16'hFFFF,
16'h088F, 16'hFFFF,
16'h0890, 16'hFFFF,
16'h0891, 16'hFFFF,
16'h0892, 16'hFFFF,
16'h0893, 16'hFFFF,
16'h0894, 16'hFFFF,
16'h0895, 16'hFFFF,
16'h0896, 16'hFFFF,
16'h0897, 16'hFFFF,
16'h0898, 16'hFFFF,
16'h0899, 16'hFFFF,
16'h089A, 16'hFFFF,
16'h089B, 16'hFFFF,
16'h089C, 16'hFFFF,
16'h089D, 16'hFFFF,
16'h089E, 16'hFFFF,
16'h089F, 16'hFFFF,
16'h08A0, 16'hFFFF,
16'h08A1, 16'hFFFF,
16'h08A2, 16'hFFFF,
16'h08A3, 16'hFFFF,
16'h08A4, 16'hFFFF,
16'h08A5, 16'hFFFF,
16'h08A6, 16'hFFFF,
16'h08A7, 16'hFFFF,
16'h08A8, 16'hFFFF,
16'h08A9, 16'hFFFF,
16'h08AA, 16'hFFFF,
16'h08AB, 16'hFFFF,
16'h08AC, 16'hFFFF,
16'h08AD, 16'hFFFF,
16'h08AE, 16'hFFFF,
16'h08AF, 16'hFFFF,
16'h08B0, 16'hFFFF,
16'h08B1, 16'hFFFF,
16'h08B2, 16'hFFFF,
16'h08B3, 16'hFFFF,
16'h08B4, 16'hFFFF,
16'h08B5, 16'hFFFF,
16'h08B6, 16'hFFFF,
16'h08B7, 16'hFFFF,
16'h08B8, 16'hFFFF,
16'h08B9, 16'hFFFF,
16'h08BA, 16'hFFFF,
16'h08BB, 16'hFFFF,
16'h08BC, 16'hFFFF,
16'h08BD, 16'hFFFF,
16'h08BE, 16'hFFFF,
16'h08BF, 16'hFFFF,
16'h08C0, 16'hFFFF,
16'h08C1, 16'hFFFF,
16'h08C2, 16'hFFFF,
16'h08C3, 16'hFFFF,
16'h08C4, 16'hFFFF,
16'h08C5, 16'hFFFF,
16'h08C6, 16'hFFFF,
16'h08C7, 16'hFFFF,
16'h08C8, 16'hFFFF,
16'h08C9, 16'hFFFF,
16'h08CA, 16'hFFFF,
16'h08CB, 16'hFFFF,
16'h08CC, 16'hFFFF,
16'h08CD, 16'hFFFF,
16'h08CE, 16'hFFFF,
16'h08CF, 16'hFFFF,
16'h08D0, 16'hFFFF,
16'h08D1, 16'hFFFF,
16'h08D2, 16'hFFFF,
16'h08D3, 16'hFFFF,
16'h08D4, 16'hFFFF,
16'h08D5, 16'hFFFF,
16'h08D6, 16'hFFFF,
16'h08D7, 16'hFFFF,
16'h08D8, 16'hFFFF,
16'h08D9, 16'hFFFF,
16'h08DA, 16'hFFFF,
16'h08DB, 16'hFFFF,
16'h08DC, 16'hFFFF,
16'h08DD, 16'hFFFF,
16'h08DE, 16'hFFFF,
16'h08DF, 16'hFFFF,
16'h08E0, 16'hFFFF,
16'h08E1, 16'hFFFF,
16'h08E2, 16'hFFFF,
16'h08E3, 16'hFFFF,
16'h08E4, 16'hFFFF,
16'h08E5, 16'hFFFF,
16'h08E6, 16'hFFFF,
16'h08E7, 16'hFFFF,
16'h08E8, 16'hFFFF,
16'h08E9, 16'hFFFF,
16'h08EA, 16'hFFFF,
16'h08EB, 16'hFFFF,
16'h08EC, 16'hFFFF,
16'h08ED, 16'hFFFF,
16'h08EE, 16'hFFFF,
16'h08EF, 16'hFFFF,
16'h08F0, 16'hFFFF,
16'h08F1, 16'hFFFF,
16'h08F2, 16'hFFFF,
16'h08F3, 16'hFFFF,
16'h08F4, 16'hFFFF,
16'h08F5, 16'hFFFF,
16'h08F6, 16'hFFFF,
16'h08F7, 16'hFFFF,
16'h08F8, 16'hFFFF,
16'h08F9, 16'hFFFF,
16'h08FA, 16'hFFFF,
16'h08FB, 16'hFFFF,
16'h08FC, 16'hFFFF,
16'h08FD, 16'hFFFF,
16'h08FE, 16'hFFFF,
16'h08FF, 16'hFFFF,
16'h0900, 16'hFFFF,
16'h0901, 16'hFFFF,
16'h0902, 16'hFFFF,
16'h0903, 16'hFFFF,
16'h0904, 16'hFFFF,
16'h0905, 16'hFFFF,
16'h0906, 16'hFFFF,
16'h0907, 16'hFFFF,
16'h0908, 16'hFFFF,
16'h0909, 16'hFFFF,
16'h090A, 16'hFFFF,
16'h090B, 16'hFFFF,
16'h090C, 16'hFFFF,
16'h090D, 16'hFFFF,
16'h090E, 16'hFFFF,
16'h090F, 16'hFFFF,
16'h0910, 16'hFFFF,
16'h0911, 16'hFFFF,
16'h0912, 16'hFFFF,
16'h0913, 16'hFFFF,
16'h0914, 16'hFFFF,
16'h0915, 16'hFFFF,
16'h0916, 16'hFFFF,
16'h0917, 16'hFFFF,
16'h0918, 16'hFFFF,
16'h0919, 16'hFFFF,
16'h091A, 16'hFFFF,
16'h091B, 16'hFFFF,
16'h091C, 16'hFFFF,
16'h091D, 16'hFFFF,
16'h091E, 16'hFFFF,
16'h091F, 16'hFFFF,
16'h0920, 16'hFFFF,
16'h0921, 16'hFFFF,
16'h0922, 16'hFFFF,
16'h0923, 16'hFFFF,
16'h0924, 16'hFFFF,
16'h0925, 16'hFFFF,
16'h0926, 16'hFFFF,
16'h0927, 16'hFFFF,
16'h0928, 16'hFFFF,
16'h0929, 16'hFFFF,
16'h092A, 16'hFFFF,
16'h092B, 16'hFFFF,
16'h092C, 16'hFFFF,
16'h092D, 16'hFFFF,
16'h092E, 16'hFFFF,
16'h092F, 16'hFFFF,
16'h0930, 16'hFFFF,
16'h0931, 16'hFFFF,
16'h0932, 16'hFFFF,
16'h0933, 16'hFFFF,
16'h0934, 16'hFFFF,
16'h0935, 16'hFFFF,
16'h0936, 16'hFFFF,
16'h0937, 16'hFFFF,
16'h0938, 16'hFFFF,
16'h0939, 16'hFFFF,
16'h093A, 16'hFFFF,
16'h093B, 16'hFFFF,
16'h093C, 16'hFFFF,
16'h093D, 16'hFFFF,
16'h093E, 16'hFFFF,
16'h093F, 16'hFFFF,
16'h0940, 16'hFFFF,
16'h0941, 16'hFFFF,
16'h0942, 16'hFFFF,
16'h0943, 16'hFFFF,
16'h0944, 16'hFFFF,
16'h0945, 16'hFFFF,
16'h0946, 16'hFFFF,
16'h0947, 16'hFFFF,
16'h0948, 16'hFFFF,
16'h0949, 16'hFFFF,
16'h094A, 16'hFFFF,
16'h094B, 16'hFFFF,
16'h094C, 16'hFFFF,
16'h094D, 16'hFFFF,
16'h094E, 16'hFFFF,
16'h094F, 16'hFFFF,
16'h0950, 16'hFFFF,
16'h0951, 16'hFFFF,
16'h0952, 16'hFFFF,
16'h0953, 16'hFFFF,
16'h0954, 16'hFFFF,
16'h0955, 16'hFFFF,
16'h0956, 16'hFFFF,
16'h0957, 16'hFFFF,
16'h0958, 16'hFFFF,
16'h0959, 16'hFFFF,
16'h095A, 16'hFFFF,
16'h095B, 16'hFFFF,
16'h095C, 16'hFFFF,
16'h095D, 16'hFFFF,
16'h095E, 16'hFFFF,
16'h095F, 16'hFFFF,
16'h0960, 16'hFFFF,
16'h0961, 16'hFFFF,
16'h0962, 16'hFFFF,
16'h0963, 16'hFFFF,
16'h0964, 16'hFFFF,
16'h0965, 16'hFFFF,
16'h0966, 16'hFFFF,
16'h0967, 16'hFFFF,
16'h0968, 16'hFFFF,
16'h0969, 16'hFFFF,
16'h096A, 16'hFFFF,
16'h096B, 16'hFFFF,
16'h096C, 16'hFFFF,
16'h096D, 16'hFFFF,
16'h096E, 16'hFFFF,
16'h096F, 16'hFFFF,
16'h0970, 16'hFFFF,
16'h0971, 16'hFFFF,
16'h0972, 16'hFFFF,
16'h0973, 16'hFFFF,
16'h0974, 16'hFFFF,
16'h0975, 16'hFFFF,
16'h0976, 16'hFFFF,
16'h0977, 16'hFFFF,
16'h0978, 16'hFFFF,
16'h0979, 16'hFFFF,
16'h097A, 16'hFFFF,
16'h097B, 16'hFFFF,
16'h097C, 16'hFFFF,
16'h097D, 16'hFFFF,
16'h097E, 16'hFFFF,
16'h097F, 16'hFFFF,
16'h0980, 16'hFFFF,
16'h0981, 16'hFFFF,
16'h0982, 16'hFFFF,
16'h0983, 16'hFFFF,
16'h0984, 16'hFFFF,
16'h0985, 16'hFFFF,
16'h0986, 16'hFFFF,
16'h0987, 16'hFFFF,
16'h0988, 16'hFFFF,
16'h0989, 16'hFFFF,
16'h098A, 16'hFFFF,
16'h098B, 16'hFFFF,
16'h098C, 16'hFFFF,
16'h098D, 16'hFFFF,
16'h098E, 16'hFFFF,
16'h098F, 16'hFFFF,
16'h0990, 16'hFFFF,
16'h0991, 16'hFFFF,
16'h0992, 16'hFFFF,
16'h0993, 16'hFFFF,
16'h0994, 16'hFFFF,
16'h0995, 16'hFFFF,
16'h0996, 16'hFFFF,
16'h0997, 16'hFFFF,
16'h0998, 16'hFFFF,
16'h0999, 16'hFFFF,
16'h099A, 16'hFFFF,
16'h099B, 16'hFFFF,
16'h099C, 16'hFFFF,
16'h099D, 16'hFFFF,
16'h099E, 16'hFFFF,
16'h099F, 16'hFFFF,
16'h09A0, 16'hFFFF,
16'h09A1, 16'hFFFF,
16'h09A2, 16'hFFFF,
16'h09A3, 16'hFFFF,
16'h09A4, 16'hFFFF,
16'h09A5, 16'hFFFF,
16'h09A6, 16'hFFFF,
16'h09A7, 16'hFFFF,
16'h09A8, 16'hFFFF,
16'h09A9, 16'hFFFF,
16'h09AA, 16'hFFFF,
16'h09AB, 16'hFFFF,
16'h09AC, 16'hFFFF,
16'h09AD, 16'hFFFF,
16'h09AE, 16'hFFFF,
16'h09AF, 16'hFFFF,
16'h09B0, 16'hFFFF,
16'h09B1, 16'hFFFF,
16'h09B2, 16'hFFFF,
16'h09B3, 16'hFFFF,
16'h09B4, 16'hFFFF,
16'h09B5, 16'hFFFF,
16'h09B6, 16'hFFFF,
16'h09B7, 16'hFFFF,
16'h09B8, 16'hFFFF,
16'h09B9, 16'hFFFF,
16'h09BA, 16'hFFFF,
16'h09BB, 16'hFFFF,
16'h09BC, 16'hFFFF,
16'h09BD, 16'hFFFF,
16'h09BE, 16'hFFFF,
16'h09BF, 16'hFFFF,
16'h09C0, 16'hFFFF,
16'h09C1, 16'hFFFF,
16'h09C2, 16'hFFFF,
16'h09C3, 16'hFFFF,
16'h09C4, 16'hFFFF,
16'h09C5, 16'hFFFF,
16'h09C6, 16'hFFFF,
16'h09C7, 16'hFFFF,
16'h09C8, 16'hFFFF,
16'h09C9, 16'hFFFF,
16'h09CA, 16'hFFFF,
16'h09CB, 16'hFFFF,
16'h09CC, 16'hFFFF,
16'h09CD, 16'hFFFF,
16'h09CE, 16'hFFFF,
16'h09CF, 16'hFFFF,
16'h09D0, 16'hFFFF,
16'h09D1, 16'hFFFF,
16'h09D2, 16'hFFFF,
16'h09D3, 16'hFFFF,
16'h09D4, 16'hFFFF,
16'h09D5, 16'hFFFF,
16'h09D6, 16'hFFFF,
16'h09D7, 16'hFFFF,
16'h09D8, 16'hFFFF,
16'h09D9, 16'hFFFF,
16'h09DA, 16'hFFFF,
16'h09DB, 16'hFFFF,
16'h09DC, 16'hFFFF,
16'h09DD, 16'hFFFF,
16'h09DE, 16'hFFFF,
16'h09DF, 16'hFFFF,
16'h09E0, 16'hFFFF,
16'h09E1, 16'hFFFF,
16'h09E2, 16'hFFFF,
16'h09E3, 16'hFFFF,
16'h09E4, 16'hFFFF,
16'h09E5, 16'hFFFF,
16'h09E6, 16'hFFFF,
16'h09E7, 16'hFFFF,
16'h09E8, 16'hFFFF,
16'h09E9, 16'hFFFF,
16'h09EA, 16'hFFFF,
16'h09EB, 16'hFFFF,
16'h09EC, 16'hFFFF,
16'h09ED, 16'hFFFF,
16'h09EE, 16'hFFFF,
16'h09EF, 16'hFFFF,
16'h09F0, 16'hFFFF,
16'h09F1, 16'hFFFF,
16'h09F2, 16'hFFFF,
16'h09F3, 16'hFFFF,
16'h09F4, 16'hFFFF,
16'h09F5, 16'hFFFF,
16'h09F6, 16'hFFFF,
16'h09F7, 16'hFFFF,
16'h09F8, 16'hFFFF,
16'h09F9, 16'hFFFF,
16'h09FA, 16'hFFFF,
16'h09FB, 16'hFFFF,
16'h09FC, 16'hFFFF,
16'h09FD, 16'hFFFF,
16'h09FE, 16'hFFFF,
16'h09FF, 16'hFFFF,
16'h0A00, 16'hFFFF,
16'h0A01, 16'hFFFF,
16'h0A02, 16'hFFFF,
16'h0A03, 16'hFFFF,
16'h0A04, 16'hFFFF,
16'h0A05, 16'hFFFF,
16'h0A06, 16'hFFFF,
16'h0A07, 16'hFFFF,
16'h0A08, 16'hFFFF,
16'h0A09, 16'hFFFF,
16'h0A0A, 16'hFFFF,
16'h0A0B, 16'hFFFF,
16'h0A0C, 16'hFFFF,
16'h0A0D, 16'hFFFF,
16'h0A0E, 16'hFFFF,
16'h0A0F, 16'hFFFF,
16'h0A10, 16'hFFFF,
16'h0A11, 16'hFFFF,
16'h0A12, 16'hFFFF,
16'h0A13, 16'hFFFF,
16'h0A14, 16'hFFFF,
16'h0A15, 16'hFFFF,
16'h0A16, 16'hFFFF,
16'h0A17, 16'hFFFF,
16'h0A18, 16'hFFFF,
16'h0A19, 16'hFFFF,
16'h0A1A, 16'hFFFF,
16'h0A1B, 16'hFFFF,
16'h0A1C, 16'hFFFF,
16'h0A1D, 16'hFFFF,
16'h0A1E, 16'hFFFF,
16'h0A1F, 16'hFFFF,
16'h0A20, 16'hFFFF,
16'h0A21, 16'hFFFF,
16'h0A22, 16'hFFFF,
16'h0A23, 16'hFFFF,
16'h0A24, 16'hFFFF,
16'h0A25, 16'hFFFF,
16'h0A26, 16'hFFFF,
16'h0A27, 16'hFFFF,
16'h0A28, 16'hFFFF,
16'h0A29, 16'hFFFF,
16'h0A2A, 16'hFFFF,
16'h0A2B, 16'hFFFF,
16'h0A2C, 16'hFFFF,
16'h0A2D, 16'hFFFF,
16'h0A2E, 16'hFFFF,
16'h0A2F, 16'hFFFF,
16'h0A30, 16'hFFFF,
16'h0A31, 16'hFFFF,
16'h0A32, 16'hFFFF,
16'h0A33, 16'hFFFF,
16'h0A34, 16'hFFFF,
16'h0A35, 16'hFFFF,
16'h0A36, 16'hFFFF,
16'h0A37, 16'hFFFF,
16'h0A38, 16'hFFFF,
16'h0A39, 16'hFFFF,
16'h0A3A, 16'hFFFF,
16'h0A3B, 16'hFFFF,
16'h0A3C, 16'hFFFF,
16'h0A3D, 16'hFFFF,
16'h0A3E, 16'hFFFF,
16'h0A3F, 16'hFFFF,
16'h0A40, 16'hFFFF,
16'h0A41, 16'hFFFF,
16'h0A42, 16'hFFFF,
16'h0A43, 16'hFFFF,
16'h0A44, 16'hFFFF,
16'h0A45, 16'hFFFF,
16'h0A46, 16'hFFFF,
16'h0A47, 16'hFFFF,
16'h0A48, 16'hFFFF,
16'h0A49, 16'hFFFF,
16'h0A4A, 16'hFFFF,
16'h0A4B, 16'hFFFF,
16'h0A4C, 16'hFFFF,
16'h0A4D, 16'hFFFF,
16'h0A4E, 16'hFFFF,
16'h0A4F, 16'hFFFF,
16'h0A50, 16'hFFFF,
16'h0A51, 16'hFFFF,
16'h0A52, 16'hFFFF,
16'h0A53, 16'hFFFF,
16'h0A54, 16'hFFFF,
16'h0A55, 16'hFFFF,
16'h0A56, 16'hFFFF,
16'h0A57, 16'hFFFF,
16'h0A58, 16'hFFFF,
16'h0A59, 16'hFFFF,
16'h0A5A, 16'hFFFF,
16'h0A5B, 16'hFFFF,
16'h0A5C, 16'hFFFF,
16'h0A5D, 16'hFFFF,
16'h0A5E, 16'hFFFF,
16'h0A5F, 16'hFFFF,
16'h0A60, 16'hFFFF,
16'h0A61, 16'hFFFF,
16'h0A62, 16'hFFFF,
16'h0A63, 16'hFFFF,
16'h0A64, 16'hFFFF,
16'h0A65, 16'hFFFF,
16'h0A66, 16'hFFFF,
16'h0A67, 16'hFFFF,
16'h0A68, 16'hFFFF,
16'h0A69, 16'hFFFF,
16'h0A6A, 16'hFFFF,
16'h0A6B, 16'hFFFF,
16'h0A6C, 16'hFFFF,
16'h0A6D, 16'hFFFF,
16'h0A6E, 16'hFFFF,
16'h0A6F, 16'hFFFF,
16'h0A70, 16'hFFFF,
16'h0A71, 16'hFFFF,
16'h0A72, 16'hFFFF,
16'h0A73, 16'hFFFF,
16'h0A74, 16'hFFFF,
16'h0A75, 16'hFFFF,
16'h0A76, 16'hFFFF,
16'h0A77, 16'hFFFF,
16'h0A78, 16'hFFFF,
16'h0A79, 16'hFFFF,
16'h0A7A, 16'hFFFF,
16'h0A7B, 16'hFFFF,
16'h0A7C, 16'hFFFF,
16'h0A7D, 16'hFFFF,
16'h0A7E, 16'hFFFF,
16'h0A7F, 16'hFFFF,
16'h0A80, 16'hFFFF,
16'h0A81, 16'hFFFF,
16'h0A82, 16'hFFFF,
16'h0A83, 16'hFFFF,
16'h0A84, 16'hFFFF,
16'h0A85, 16'hFFFF,
16'h0A86, 16'hFFFF,
16'h0A87, 16'hFFFF,
16'h0A88, 16'hFFFF,
16'h0A89, 16'hFFFF,
16'h0A8A, 16'hFFFF,
16'h0A8B, 16'hFFFF,
16'h0A8C, 16'hFFFF,
16'h0A8D, 16'hFFFF,
16'h0A8E, 16'hFFFF,
16'h0A8F, 16'hFFFF,
16'h0A90, 16'hFFFF,
16'h0A91, 16'hFFFF,
16'h0A92, 16'hFFFF,
16'h0A93, 16'hFFFF,
16'h0A94, 16'hFFFF,
16'h0A95, 16'hFFFF,
16'h0A96, 16'hFFFF,
16'h0A97, 16'hFFFF,
16'h0A98, 16'hFFFF,
16'h0A99, 16'hFFFF,
16'h0A9A, 16'hFFFF,
16'h0A9B, 16'hFFFF,
16'h0A9C, 16'hFFFF,
16'h0A9D, 16'hFFFF,
16'h0A9E, 16'hFFFF,
16'h0A9F, 16'hFFFF,
16'h0AA0, 16'hFFFF,
16'h0AA1, 16'hFFFF,
16'h0AA2, 16'hFFFF,
16'h0AA3, 16'hFFFF,
16'h0AA4, 16'hFFFF,
16'h0AA5, 16'hFFFF,
16'h0AA6, 16'hFFFF,
16'h0AA7, 16'hFFFF,
16'h0AA8, 16'hFFFF,
16'h0AA9, 16'hFFFF,
16'h0AAA, 16'hFFFF,
16'h0AAB, 16'hFFFF,
16'h0AAC, 16'hFFFF,
16'h0AAD, 16'hFFFF,
16'h0AAE, 16'hFFFF,
16'h0AAF, 16'hFFFF,
16'h0AB0, 16'hFFFF,
16'h0AB1, 16'hFFFF,
16'h0AB2, 16'hFFFF,
16'h0AB3, 16'hFFFF,
16'h0AB4, 16'hFFFF,
16'h0AB5, 16'hFFFF,
16'h0AB6, 16'hFFFF,
16'h0AB7, 16'hFFFF,
16'h0AB8, 16'hFFFF,
16'h0AB9, 16'hFFFF,
16'h0ABA, 16'hFFFF,
16'h0ABB, 16'hFFFF,
16'h0ABC, 16'hFFFF,
16'h0ABD, 16'hFFFF,
16'h0ABE, 16'hFFFF,
16'h0ABF, 16'hFFFF,
16'h0AC0, 16'hFFFF,
16'h0AC1, 16'hFFFF,
16'h0AC2, 16'hFFFF,
16'h0AC3, 16'hFFFF,
16'h0AC4, 16'hFFFF,
16'h0AC5, 16'hFFFF,
16'h0AC6, 16'hFFFF,
16'h0AC7, 16'hFFFF,
16'h0AC8, 16'hFFFF,
16'h0AC9, 16'hFFFF,
16'h0ACA, 16'hFFFF,
16'h0ACB, 16'hFFFF,
16'h0ACC, 16'hFFFF,
16'h0ACD, 16'hFFFF,
16'h0ACE, 16'hFFFF,
16'h0ACF, 16'hFFFF,
16'h0AD0, 16'hFFFF,
16'h0AD1, 16'hFFFF,
16'h0AD2, 16'hFFFF,
16'h0AD3, 16'hFFFF,
16'h0AD4, 16'hFFFF,
16'h0AD5, 16'hFFFF,
16'h0AD6, 16'hFFFF,
16'h0AD7, 16'hFFFF,
16'h0AD8, 16'hFFFF,
16'h0AD9, 16'hFFFF,
16'h0ADA, 16'hFFFF,
16'h0ADB, 16'hFFFF,
16'h0ADC, 16'hFFFF,
16'h0ADD, 16'hFFFF,
16'h0ADE, 16'hFFFF,
16'h0ADF, 16'hFFFF,
16'h0AE0, 16'hFFFF,
16'h0AE1, 16'hFFFF,
16'h0AE2, 16'hFFFF,
16'h0AE3, 16'hFFFF,
16'h0AE4, 16'hFFFF,
16'h0AE5, 16'hFFFF,
16'h0AE6, 16'hFFFF,
16'h0AE7, 16'hFFFF,
16'h0AE8, 16'hFFFF,
16'h0AE9, 16'hFFFF,
16'h0AEA, 16'hFFFF,
16'h0AEB, 16'hFFFF,
16'h0AEC, 16'hFFFF,
16'h0AED, 16'hFFFF,
16'h0AEE, 16'hFFFF,
16'h0AEF, 16'hFFFF,
16'h0AF0, 16'hFFFF,
16'h0AF1, 16'hFFFF,
16'h0AF2, 16'hFFFF,
16'h0AF3, 16'hFFFF,
16'h0AF4, 16'hFFFF,
16'h0AF5, 16'hFFFF,
16'h0AF6, 16'hFFFF,
16'h0AF7, 16'hFFFF,
16'h0AF8, 16'hFFFF,
16'h0AF9, 16'hFFFF,
16'h0AFA, 16'hFFFF,
16'h0AFB, 16'hFFFF,
16'h0AFC, 16'hFFFF,
16'h0AFD, 16'hFFFF,
16'h0AFE, 16'hFFFF,
16'h0AFF, 16'hFFFF,
16'h0B00, 16'hFFFF,
16'h0B01, 16'hFFFF,
16'h0B02, 16'hFFFF,
16'h0B03, 16'hFFFF,
16'h0B04, 16'hFFFF,
16'h0B05, 16'hFFFF,
16'h0B06, 16'hFFFF,
16'h0B07, 16'hFFFF,
16'h0B08, 16'hFFFF,
16'h0B09, 16'hFFFF,
16'h0B0A, 16'hFFFF,
16'h0B0B, 16'hFFFF,
16'h0B0C, 16'hFFFF,
16'h0B0D, 16'hFFFF,
16'h0B0E, 16'hFFFF,
16'h0B0F, 16'hFFFF,
16'h0B10, 16'hFFFF,
16'h0B11, 16'hFFFF,
16'h0B12, 16'hFFFF,
16'h0B13, 16'hFFFF,
16'h0B14, 16'hFFFF,
16'h0B15, 16'hFFFF,
16'h0B16, 16'hFFFF,
16'h0B17, 16'hFFFF,
16'h0B18, 16'hFFFF,
16'h0B19, 16'hFFFF,
16'h0B1A, 16'hFFFF,
16'h0B1B, 16'hFFFF,
16'h0B1C, 16'hFFFF,
16'h0B1D, 16'hFFFF,
16'h0B1E, 16'hFFFF,
16'h0B1F, 16'hFFFF,
16'h0B20, 16'hFFFF,
16'h0B21, 16'hFFFF,
16'h0B22, 16'hFFFF,
16'h0B23, 16'hFFFF,
16'h0B24, 16'hFFFF,
16'h0B25, 16'hFFFF,
16'h0B26, 16'hFFFF,
16'h0B27, 16'hFFFF,
16'h0B28, 16'hFFFF,
16'h0B29, 16'hFFFF,
16'h0B2A, 16'hFFFF,
16'h0B2B, 16'hFFFF,
16'h0B2C, 16'hFFFF,
16'h0B2D, 16'hFFFF,
16'h0B2E, 16'hFFFF,
16'h0B2F, 16'hFFFF,
16'h0B30, 16'hFFFF,
16'h0B31, 16'hFFFF,
16'h0B32, 16'hFFFF,
16'h0B33, 16'hFFFF,
16'h0B34, 16'hFFFF,
16'h0B35, 16'hFFFF,
16'h0B36, 16'hFFFF,
16'h0B37, 16'hFFFF,
16'h0B38, 16'hFFFF,
16'h0B39, 16'hFFFF,
16'h0B3A, 16'hFFFF,
16'h0B3B, 16'hFFFF,
16'h0B3C, 16'hFFFF,
16'h0B3D, 16'hFFFF,
16'h0B3E, 16'hFFFF,
16'h0B3F, 16'hFFFF,
16'h0B40, 16'hFFFF,
16'h0B41, 16'hFFFF,
16'h0B42, 16'hFFFF,
16'h0B43, 16'hFFFF,
16'h0B44, 16'hFFFF,
16'h0B45, 16'hFFFF,
16'h0B46, 16'hFFFF,
16'h0B47, 16'hFFFF,
16'h0B48, 16'hFFFF,
16'h0B49, 16'hFFFF,
16'h0B4A, 16'hFFFF,
16'h0B4B, 16'hFFFF,
16'h0B4C, 16'hFFFF,
16'h0B4D, 16'hFFFF,
16'h0B4E, 16'hFFFF,
16'h0B4F, 16'hFFFF,
16'h0B50, 16'hFFFF,
16'h0B51, 16'hFFFF,
16'h0B52, 16'hFFFF,
16'h0B53, 16'hFFFF,
16'h0B54, 16'hFFFF,
16'h0B55, 16'hFFFF,
16'h0B56, 16'hFFFF,
16'h0B57, 16'hFFFF,
16'h0B58, 16'hFFFF,
16'h0B59, 16'hFFFF,
16'h0B5A, 16'hFFFF,
16'h0B5B, 16'hFFFF,
16'h0B5C, 16'hFFFF,
16'h0B5D, 16'hFFFF,
16'h0B5E, 16'hFFFF,
16'h0B5F, 16'hFFFF,
16'h0B60, 16'hFFFF,
16'h0B61, 16'hFFFF,
16'h0B62, 16'hFFFF,
16'h0B63, 16'hFFFF,
16'h0B64, 16'hFFFF,
16'h0B65, 16'hFFFF,
16'h0B66, 16'hFFFF,
16'h0B67, 16'hFFFF,
16'h0B68, 16'hFFFF,
16'h0B69, 16'hFFFF,
16'h0B6A, 16'hFFFF,
16'h0B6B, 16'hFFFF,
16'h0B6C, 16'hFFFF,
16'h0B6D, 16'hFFFF,
16'h0B6E, 16'hFFFF,
16'h0B6F, 16'hFFFF,
16'h0B70, 16'hFFFF,
16'h0B71, 16'hFFFF,
16'h0B72, 16'hFFFF,
16'h0B73, 16'hFFFF,
16'h0B74, 16'hFFFF,
16'h0B75, 16'hFFFF,
16'h0B76, 16'hFFFF,
16'h0B77, 16'hFFFF,
16'h0B78, 16'hFFFF,
16'h0B79, 16'hFFFF,
16'h0B7A, 16'hFFFF,
16'h0B7B, 16'hFFFF,
16'h0B7C, 16'hFFFF,
16'h0B7D, 16'hFFFF,
16'h0B7E, 16'hFFFF,
16'h0B7F, 16'hFFFF,
16'h0B80, 16'hFFFF,
16'h0B81, 16'hFFFF,
16'h0B82, 16'hFFFF,
16'h0B83, 16'hFFFF,
16'h0B84, 16'hFFFF,
16'h0B85, 16'hFFFF,
16'h0B86, 16'hFFFF,
16'h0B87, 16'hFFFF,
16'h0B88, 16'hFFFF,
16'h0B89, 16'hFFFF,
16'h0B8A, 16'hFFFF,
16'h0B8B, 16'hFFFF,
16'h0B8C, 16'hFFFF,
16'h0B8D, 16'hFFFF,
16'h0B8E, 16'hFFFF,
16'h0B8F, 16'hFFFF,
16'h0B90, 16'hFFFF,
16'h0B91, 16'hFFFF,
16'h0B92, 16'hFFFF,
16'h0B93, 16'hFFFF,
16'h0B94, 16'hFFFF,
16'h0B95, 16'hFFFF,
16'h0B96, 16'hFFFF,
16'h0B97, 16'hFFFF,
16'h0B98, 16'hFFFF,
16'h0B99, 16'hFFFF,
16'h0B9A, 16'hFFFF,
16'h0B9B, 16'hFFFF,
16'h0B9C, 16'hFFFF,
16'h0B9D, 16'hFFFF,
16'h0B9E, 16'hFFFF,
16'h0B9F, 16'hFFFF,
16'h0BA0, 16'hFFFF,
16'h0BA1, 16'hFFFF,
16'h0BA2, 16'hFFFF,
16'h0BA3, 16'hFFFF,
16'h0BA4, 16'hFFFF,
16'h0BA5, 16'hFFFF,
16'h0BA6, 16'hFFFF,
16'h0BA7, 16'hFFFF,
16'h0BA8, 16'hFFFF,
16'h0BA9, 16'hFFFF,
16'h0BAA, 16'hFFFF,
16'h0BAB, 16'hFFFF,
16'h0BAC, 16'hFFFF,
16'h0BAD, 16'hFFFF,
16'h0BAE, 16'hFFFF,
16'h0BAF, 16'hFFFF,
16'h0BB0, 16'hFFFF,
16'h0BB1, 16'hFFFF,
16'h0BB2, 16'hFFFF,
16'h0BB3, 16'hFFFF,
16'h0BB4, 16'hFFFF,
16'h0BB5, 16'hFFFF,
16'h0BB6, 16'hFFFF,
16'h0BB7, 16'hFFFF,
16'h0BB8, 16'hFFFF,
16'h0BB9, 16'hFFFF,
16'h0BBA, 16'hFFFF,
16'h0BBB, 16'hFFFF,
16'h0BBC, 16'hFFFF,
16'h0BBD, 16'hFFFF,
16'h0BBE, 16'hFFFF,
16'h0BBF, 16'hFFFF,
16'h0BC0, 16'hFFFF,
16'h0BC1, 16'hFFFF,
16'h0BC2, 16'hFFFF,
16'h0BC3, 16'hFFFF,
16'h0BC4, 16'hFFFF,
16'h0BC5, 16'hFFFF,
16'h0BC6, 16'hFFFF,
16'h0BC7, 16'hFFFF,
16'h0BC8, 16'hFFFF,
16'h0BC9, 16'hFFFF,
16'h0BCA, 16'hFFFF,
16'h0BCB, 16'hFFFF,
16'h0BCC, 16'hFFFF,
16'h0BCD, 16'hFFFF,
16'h0BCE, 16'hFFFF,
16'h0BCF, 16'hFFFF,
16'h0BD0, 16'hFFFF,
16'h0BD1, 16'hFFFF,
16'h0BD2, 16'hFFFF,
16'h0BD3, 16'hFFFF,
16'h0BD4, 16'hFFFF,
16'h0BD5, 16'hFFFF,
16'h0BD6, 16'hFFFF,
16'h0BD7, 16'hFFFF,
16'h0BD8, 16'hFFFF,
16'h0BD9, 16'hFFFF,
16'h0BDA, 16'hFFFF,
16'h0BDB, 16'hFFFF,
16'h0BDC, 16'hFFFF,
16'h0BDD, 16'hFFFF,
16'h0BDE, 16'hFFFF,
16'h0BDF, 16'hFFFF,
16'h0BE0, 16'hFFFF,
16'h0BE1, 16'hFFFF,
16'h0BE2, 16'hFFFF,
16'h0BE3, 16'hFFFF,
16'h0BE4, 16'hFFFF,
16'h0BE5, 16'hFFFF,
16'h0BE6, 16'hFFFF,
16'h0BE7, 16'hFFFF,
16'h0BE8, 16'hFFFF,
16'h0BE9, 16'hFFFF,
16'h0BEA, 16'hFFFF,
16'h0BEB, 16'hFFFF,
16'h0BEC, 16'hFFFF,
16'h0BED, 16'hFFFF,
16'h0BEE, 16'hFFFF,
16'h0BEF, 16'hFFFF,
16'h0BF0, 16'hFFFF,
16'h0BF1, 16'hFFFF,
16'h0BF2, 16'hFFFF,
16'h0BF3, 16'hFFFF,
16'h0BF4, 16'hFFFF,
16'h0BF5, 16'hFFFF,
16'h0BF6, 16'hFFFF,
16'h0BF7, 16'hFFFF,
16'h0BF8, 16'hFFFF,
16'h0BF9, 16'hFFFF,
16'h0BFA, 16'hFFFF,
16'h0BFB, 16'hFFFF,
16'h0BFC, 16'hFFFF,
16'h0BFD, 16'hFFFF,
16'h0BFE, 16'hFFFF,
16'h0BFF, 16'hFFFF,
16'h0C00, 16'hFFFF,
16'h0C01, 16'hFFFF,
16'h0C02, 16'hFFFF,
16'h0C03, 16'hFFFF,
16'h0C04, 16'hFFFF,
16'h0C05, 16'hFFFF,
16'h0C06, 16'hFFFF,
16'h0C07, 16'hFFFF,
16'h0C08, 16'hFFFF,
16'h0C09, 16'hFFFF,
16'h0C0A, 16'hFFFF,
16'h0C0B, 16'hFFFF,
16'h0C0C, 16'hFFFF,
16'h0C0D, 16'hFFFF,
16'h0C0E, 16'hFFFF,
16'h0C0F, 16'hFFFF,
16'h0C10, 16'hFFFF,
16'h0C11, 16'hFFFF,
16'h0C12, 16'hFFFF,
16'h0C13, 16'hFFFF,
16'h0C14, 16'hFFFF,
16'h0C15, 16'hFFFF,
16'h0C16, 16'hFFFF,
16'h0C17, 16'hFFFF,
16'h0C18, 16'hFFFF,
16'h0C19, 16'hFFFF,
16'h0C1A, 16'hFFFF,
16'h0C1B, 16'hFFFF,
16'h0C1C, 16'hFFFF,
16'h0C1D, 16'hFFFF,
16'h0C1E, 16'hFFFF,
16'h0C1F, 16'hFFFF,
16'h0C20, 16'hFFFF,
16'h0C21, 16'hFFFF,
16'h0C22, 16'hFFFF,
16'h0C23, 16'hFFFF,
16'h0C24, 16'hFFFF,
16'h0C25, 16'hFFFF,
16'h0C26, 16'hFFFF,
16'h0C27, 16'hFFFF,
16'h0C28, 16'hFFFF,
16'h0C29, 16'hFFFF,
16'h0C2A, 16'hFFFF,
16'h0C2B, 16'hFFFF,
16'h0C2C, 16'hFFFF,
16'h0C2D, 16'hFFFF,
16'h0C2E, 16'hFFFF,
16'h0C2F, 16'hFFFF,
16'h0C30, 16'hFFFF,
16'h0C31, 16'hFFFF,
16'h0C32, 16'hFFFF,
16'h0C33, 16'hFFFF,
16'h0C34, 16'hFFFF,
16'h0C35, 16'hFFFF,
16'h0C36, 16'hFFFF,
16'h0C37, 16'hFFFF,
16'h0C38, 16'hFFFF,
16'h0C39, 16'hFFFF,
16'h0C3A, 16'hFFFF,
16'h0C3B, 16'hFFFF,
16'h0C3C, 16'hFFFF,
16'h0C3D, 16'hFFFF,
16'h0C3E, 16'hFFFF,
16'h0C3F, 16'hFFFF,
16'h0C40, 16'hFFFF,
16'h0C41, 16'hFFFF,
16'h0C42, 16'hFFFF,
16'h0C43, 16'hFFFF,
16'h0C44, 16'hFFFF,
16'h0C45, 16'hFFFF,
16'h0C46, 16'hFFFF,
16'h0C47, 16'hFFFF,
16'h0C48, 16'hFFFF,
16'h0C49, 16'hFFFF,
16'h0C4A, 16'hFFFF,
16'h0C4B, 16'hFFFF,
16'h0C4C, 16'hFFFF,
16'h0C4D, 16'hFFFF,
16'h0C4E, 16'hFFFF,
16'h0C4F, 16'hFFFF,
16'h0C50, 16'hFFFF,
16'h0C51, 16'hFFFF,
16'h0C52, 16'hFFFF,
16'h0C53, 16'hFFFF,
16'h0C54, 16'hFFFF,
16'h0C55, 16'hFFFF,
16'h0C56, 16'hFFFF,
16'h0C57, 16'hFFFF,
16'h0C58, 16'hFFFF,
16'h0C59, 16'hFFFF,
16'h0C5A, 16'hFFFF,
16'h0C5B, 16'hFFFF,
16'h0C5C, 16'hFFFF,
16'h0C5D, 16'hFFFF,
16'h0C5E, 16'hFFFF,
16'h0C5F, 16'hFFFF,
16'h0C60, 16'hFFFF,
16'h0C61, 16'hFFFF,
16'h0C62, 16'hFFFF,
16'h0C63, 16'hFFFF,
16'h0C64, 16'hFFFF,
16'h0C65, 16'hFFFF,
16'h0C66, 16'hFFFF,
16'h0C67, 16'hFFFF,
16'h0C68, 16'hFFFF,
16'h0C69, 16'hFFFF,
16'h0C6A, 16'hFFFF,
16'h0C6B, 16'hFFFF,
16'h0C6C, 16'hFFFF,
16'h0C6D, 16'hFFFF,
16'h0C6E, 16'hFFFF,
16'h0C6F, 16'hFFFF,
16'h0C70, 16'hFFFF,
16'h0C71, 16'hFFFF,
16'h0C72, 16'hFFFF,
16'h0C73, 16'hFFFF,
16'h0C74, 16'hFFFF,
16'h0C75, 16'hFFFF,
16'h0C76, 16'hFFFF,
16'h0C77, 16'hFFFF,
16'h0C78, 16'hFFFF,
16'h0C79, 16'hFFFF,
16'h0C7A, 16'hFFFF,
16'h0C7B, 16'hFFFF,
16'h0C7C, 16'hFFFF,
16'h0C7D, 16'hFFFF,
16'h0C7E, 16'hFFFF,
16'h0C7F, 16'hFFFF,
16'h0C80, 16'hFFFF,
16'h0C81, 16'hFFFF,
16'h0C82, 16'hFFFF,
16'h0C83, 16'hFFFF,
16'h0C84, 16'hFFFF,
16'h0C85, 16'hFFFF,
16'h0C86, 16'hFFFF,
16'h0C87, 16'hFFFF,
16'h0C88, 16'hFFFF,
16'h0C89, 16'hFFFF,
16'h0C8A, 16'hFFFF,
16'h0C8B, 16'hFFFF,
16'h0C8C, 16'hFFFF,
16'h0C8D, 16'hFFFF,
16'h0C8E, 16'hFFFF,
16'h0C8F, 16'hFFFF,
16'h0C90, 16'hFFFF,
16'h0C91, 16'hFFFF,
16'h0C92, 16'hFFFF,
16'h0C93, 16'hFFFF,
16'h0C94, 16'hFFFF,
16'h0C95, 16'hFFFF,
16'h0C96, 16'hFFFF,
16'h0C97, 16'hFFFF,
16'h0C98, 16'hFFFF,
16'h0C99, 16'hFFFF,
16'h0C9A, 16'hFFFF,
16'h0C9B, 16'hFFFF,
16'h0C9C, 16'hFFFF,
16'h0C9D, 16'hFFFF,
16'h0C9E, 16'hFFFF,
16'h0C9F, 16'hFFFF,
16'h0CA0, 16'hFFFF,
16'h0CA1, 16'hFFFF,
16'h0CA2, 16'hFFFF,
16'h0CA3, 16'hFFFF,
16'h0CA4, 16'hFFFF,
16'h0CA5, 16'hFFFF,
16'h0CA6, 16'hFFFF,
16'h0CA7, 16'hFFFF,
16'h0CA8, 16'hFFFF,
16'h0CA9, 16'hFFFF,
16'h0CAA, 16'hFFFF,
16'h0CAB, 16'hFFFF,
16'h0CAC, 16'hFFFF,
16'h0CAD, 16'hFFFF,
16'h0CAE, 16'hFFFF,
16'h0CAF, 16'hFFFF,
16'h0CB0, 16'hFFFF,
16'h0CB1, 16'hFFFF,
16'h0CB2, 16'hFFFF,
16'h0CB3, 16'hFFFF,
16'h0CB4, 16'hFFFF,
16'h0CB5, 16'hFFFF,
16'h0CB6, 16'hFFFF,
16'h0CB7, 16'hFFFF,
16'h0CB8, 16'hFFFF,
16'h0CB9, 16'hFFFF,
16'h0CBA, 16'hFFFF,
16'h0CBB, 16'hFFFF,
16'h0CBC, 16'hFFFF,
16'h0CBD, 16'hFFFF,
16'h0CBE, 16'hFFFF,
16'h0CBF, 16'hFFFF,
16'h0CC0, 16'hFFFF,
16'h0CC1, 16'hFFFF,
16'h0CC2, 16'hFFFF,
16'h0CC3, 16'hFFFF,
16'h0CC4, 16'hFFFF,
16'h0CC5, 16'hFFFF,
16'h0CC6, 16'hFFFF,
16'h0CC7, 16'hFFFF,
16'h0CC8, 16'hFFFF,
16'h0CC9, 16'hFFFF,
16'h0CCA, 16'hFFFF,
16'h0CCB, 16'hFFFF,
16'h0CCC, 16'hFFFF,
16'h0CCD, 16'hFFFF,
16'h0CCE, 16'hFFFF,
16'h0CCF, 16'hFFFF,
16'h0CD0, 16'hFFFF,
16'h0CD1, 16'hFFFF,
16'h0CD2, 16'hFFFF,
16'h0CD3, 16'hFFFF,
16'h0CD4, 16'hFFFF,
16'h0CD5, 16'hFFFF,
16'h0CD6, 16'hFFFF,
16'h0CD7, 16'hFFFF,
16'h0CD8, 16'hFFFF,
16'h0CD9, 16'hFFFF,
16'h0CDA, 16'hFFFF,
16'h0CDB, 16'hFFFF,
16'h0CDC, 16'hFFFF,
16'h0CDD, 16'hFFFF,
16'h0CDE, 16'hFFFF,
16'h0CDF, 16'hFFFF,
16'h0CE0, 16'hFFFF,
16'h0CE1, 16'hFFFF,
16'h0CE2, 16'hFFFF,
16'h0CE3, 16'hFFFF,
16'h0CE4, 16'hFFFF,
16'h0CE5, 16'hFFFF,
16'h0CE6, 16'hFFFF,
16'h0CE7, 16'hFFFF,
16'h0CE8, 16'hFFFF,
16'h0CE9, 16'hFFFF,
16'h0CEA, 16'hFFFF,
16'h0CEB, 16'hFFFF,
16'h0CEC, 16'hFFFF,
16'h0CED, 16'hFFFF,
16'h0CEE, 16'hFFFF,
16'h0CEF, 16'hFFFF,
16'h0CF0, 16'hFFFF,
16'h0CF1, 16'hFFFF,
16'h0CF2, 16'hFFFF,
16'h0CF3, 16'hFFFF,
16'h0CF4, 16'hFFFF,
16'h0CF5, 16'hFFFF,
16'h0CF6, 16'hFFFF,
16'h0CF7, 16'hFFFF,
16'h0CF8, 16'hFFFF,
16'h0CF9, 16'hFFFF,
16'h0CFA, 16'hFFFF,
16'h0CFB, 16'hFFFF,
16'h0CFC, 16'hFFFF,
16'h0CFD, 16'hFFFF,
16'h0CFE, 16'hFFFF,
16'h0CFF, 16'hFFFF,
16'h0D00, 16'hFFFF,
16'h0D01, 16'hFFFF,
16'h0D02, 16'hFFFF,
16'h0D03, 16'hFFFF,
16'h0D04, 16'hFFFF,
16'h0D05, 16'hFFFF,
16'h0D06, 16'hFFFF,
16'h0D07, 16'hFFFF,
16'h0D08, 16'hFFFF,
16'h0D09, 16'hFFFF,
16'h0D0A, 16'hFFFF,
16'h0D0B, 16'hFFFF,
16'h0D0C, 16'hFFFF,
16'h0D0D, 16'hFFFF,
16'h0D0E, 16'hFFFF,
16'h0D0F, 16'hFFFF,
16'h0D10, 16'hFFFF,
16'h0D11, 16'hFFFF,
16'h0D12, 16'hFFFF,
16'h0D13, 16'hFFFF,
16'h0D14, 16'hFFFF,
16'h0D15, 16'hFFFF,
16'h0D16, 16'hFFFF,
16'h0D17, 16'hFFFF,
16'h0D18, 16'hFFFF,
16'h0D19, 16'hFFFF,
16'h0D1A, 16'hFFFF,
16'h0D1B, 16'hFFFF,
16'h0D1C, 16'hFFFF,
16'h0D1D, 16'hFFFF,
16'h0D1E, 16'hFFFF,
16'h0D1F, 16'hFFFF,
16'h0D20, 16'hFFFF,
16'h0D21, 16'hFFFF,
16'h0D22, 16'hFFFF,
16'h0D23, 16'hFFFF,
16'h0D24, 16'hFFFF,
16'h0D25, 16'hFFFF,
16'h0D26, 16'hFFFF,
16'h0D27, 16'hFFFF,
16'h0D28, 16'hFFFF,
16'h0D29, 16'hFFFF,
16'h0D2A, 16'hFFFF,
16'h0D2B, 16'hFFFF,
16'h0D2C, 16'hFFFF,
16'h0D2D, 16'hFFFF,
16'h0D2E, 16'hFFFF,
16'h0D2F, 16'hFFFF,
16'h0D30, 16'hFFFF,
16'h0D31, 16'hFFFF,
16'h0D32, 16'hFFFF,
16'h0D33, 16'hFFFF,
16'h0D34, 16'hFFFF,
16'h0D35, 16'hFFFF,
16'h0D36, 16'hFFFF,
16'h0D37, 16'hFFFF,
16'h0D38, 16'hFFFF,
16'h0D39, 16'hFFFF,
16'h0D3A, 16'hFFFF,
16'h0D3B, 16'hFFFF,
16'h0D3C, 16'hFFFF,
16'h0D3D, 16'hFFFF,
16'h0D3E, 16'hFFFF,
16'h0D3F, 16'hFFFF,
16'h0D40, 16'hFFFF,
16'h0D41, 16'hFFFF,
16'h0D42, 16'hFFFF,
16'h0D43, 16'hFFFF,
16'h0D44, 16'hFFFF,
16'h0D45, 16'hFFFF,
16'h0D46, 16'hFFFF,
16'h0D47, 16'hFFFF,
16'h0D48, 16'hFFFF,
16'h0D49, 16'hFFFF,
16'h0D4A, 16'hFFFF,
16'h0D4B, 16'hFFFF,
16'h0D4C, 16'hFFFF,
16'h0D4D, 16'hFFFF,
16'h0D4E, 16'hFFFF,
16'h0D4F, 16'hFFFF,
16'h0D50, 16'hFFFF,
16'h0D51, 16'hFFFF,
16'h0D52, 16'hFFFF,
16'h0D53, 16'hFFFF,
16'h0D54, 16'hFFFF,
16'h0D55, 16'hFFFF,
16'h0D56, 16'hFFFF,
16'h0D57, 16'hFFFF,
16'h0D58, 16'hFFFF,
16'h0D59, 16'hFFFF,
16'h0D5A, 16'hFFFF,
16'h0D5B, 16'hFFFF,
16'h0D5C, 16'hFFFF,
16'h0D5D, 16'hFFFF,
16'h0D5E, 16'hFFFF,
16'h0D5F, 16'hFFFF,
16'h0D60, 16'hFFFF,
16'h0D61, 16'hFFFF,
16'h0D62, 16'hFFFF,
16'h0D63, 16'hFFFF,
16'h0D64, 16'hFFFF,
16'h0D65, 16'hFFFF,
16'h0D66, 16'hFFFF,
16'h0D67, 16'hFFFF,
16'h0D68, 16'hFFFF,
16'h0D69, 16'hFFFF,
16'h0D6A, 16'hFFFF,
16'h0D6B, 16'hFFFF,
16'h0D6C, 16'hFFFF,
16'h0D6D, 16'hFFFF,
16'h0D6E, 16'hFFFF,
16'h0D6F, 16'hFFFF,
16'h0D70, 16'hFFFF,
16'h0D71, 16'hFFFF,
16'h0D72, 16'hFFFF,
16'h0D73, 16'hFFFF,
16'h0D74, 16'hFFFF,
16'h0D75, 16'hFFFF,
16'h0D76, 16'hFFFF,
16'h0D77, 16'hFFFF,
16'h0D78, 16'hFFFF,
16'h0D79, 16'hFFFF,
16'h0D7A, 16'hFFFF,
16'h0D7B, 16'hFFFF,
16'h0D7C, 16'hFFFF,
16'h0D7D, 16'hFFFF,
16'h0D7E, 16'hFFFF,
16'h0D7F, 16'hFFFF,
16'h0D80, 16'hFFFF,
16'h0D81, 16'hFFFF,
16'h0D82, 16'hFFFF,
16'h0D83, 16'hFFFF,
16'h0D84, 16'hFFFF,
16'h0D85, 16'hFFFF,
16'h0D86, 16'hFFFF,
16'h0D87, 16'hFFFF,
16'h0D88, 16'hFFFF,
16'h0D89, 16'hFFFF,
16'h0D8A, 16'hFFFF,
16'h0D8B, 16'hFFFF,
16'h0D8C, 16'hFFFF,
16'h0D8D, 16'hFFFF,
16'h0D8E, 16'hFFFF,
16'h0D8F, 16'hFFFF,
16'h0D90, 16'hFFFF,
16'h0D91, 16'hFFFF,
16'h0D92, 16'hFFFF,
16'h0D93, 16'hFFFF,
16'h0D94, 16'hFFFF,
16'h0D95, 16'hFFFF,
16'h0D96, 16'hFFFF,
16'h0D97, 16'hFFFF,
16'h0D98, 16'hFFFF,
16'h0D99, 16'hFFFF,
16'h0D9A, 16'hFFFF,
16'h0D9B, 16'hFFFF,
16'h0D9C, 16'hFFFF,
16'h0D9D, 16'hFFFF,
16'h0D9E, 16'hFFFF,
16'h0D9F, 16'hFFFF,
16'h0DA0, 16'hFFFF,
16'h0DA1, 16'hFFFF,
16'h0DA2, 16'hFFFF,
16'h0DA3, 16'hFFFF,
16'h0DA4, 16'hFFFF,
16'h0DA5, 16'hFFFF,
16'h0DA6, 16'hFFFF,
16'h0DA7, 16'hFFFF,
16'h0DA8, 16'hFFFF,
16'h0DA9, 16'hFFFF,
16'h0DAA, 16'hFFFF,
16'h0DAB, 16'hFFFF,
16'h0DAC, 16'hFFFF,
16'h0DAD, 16'hFFFF,
16'h0DAE, 16'hFFFF,
16'h0DAF, 16'hFFFF,
16'h0DB0, 16'hFFFF,
16'h0DB1, 16'hFFFF,
16'h0DB2, 16'hFFFF,
16'h0DB3, 16'hFFFF,
16'h0DB4, 16'hFFFF,
16'h0DB5, 16'hFFFF,
16'h0DB6, 16'hFFFF,
16'h0DB7, 16'hFFFF,
16'h0DB8, 16'hFFFF,
16'h0DB9, 16'hFFFF,
16'h0DBA, 16'hFFFF,
16'h0DBB, 16'hFFFF,
16'h0DBC, 16'hFFFF,
16'h0DBD, 16'hFFFF,
16'h0DBE, 16'hFFFF,
16'h0DBF, 16'hFFFF,
16'h0DC0, 16'hFFFF,
16'h0DC1, 16'hFFFF,
16'h0DC2, 16'hFFFF,
16'h0DC3, 16'hFFFF,
16'h0DC4, 16'hFFFF,
16'h0DC5, 16'hFFFF,
16'h0DC6, 16'hFFFF,
16'h0DC7, 16'hFFFF,
16'h0DC8, 16'hFFFF,
16'h0DC9, 16'hFFFF,
16'h0DCA, 16'hFFFF,
16'h0DCB, 16'hFFFF,
16'h0DCC, 16'hFFFF,
16'h0DCD, 16'hFFFF,
16'h0DCE, 16'hFFFF,
16'h0DCF, 16'hFFFF,
16'h0DD0, 16'hFFFF,
16'h0DD1, 16'hFFFF,
16'h0DD2, 16'hFFFF,
16'h0DD3, 16'hFFFF,
16'h0DD4, 16'hFFFF,
16'h0DD5, 16'hFFFF,
16'h0DD6, 16'hFFFF,
16'h0DD7, 16'hFFFF,
16'h0DD8, 16'hFFFF,
16'h0DD9, 16'hFFFF,
16'h0DDA, 16'hFFFF,
16'h0DDB, 16'hFFFF,
16'h0DDC, 16'hFFFF,
16'h0DDD, 16'hFFFF,
16'h0DDE, 16'hFFFF,
16'h0DDF, 16'hFFFF,
16'h0DE0, 16'hFFFF,
16'h0DE1, 16'hFFFF,
16'h0DE2, 16'hFFFF,
16'h0DE3, 16'hFFFF,
16'h0DE4, 16'hFFFF,
16'h0DE5, 16'hFFFF,
16'h0DE6, 16'hFFFF,
16'h0DE7, 16'hFFFF,
16'h0DE8, 16'hFFFF,
16'h0DE9, 16'hFFFF,
16'h0DEA, 16'hFFFF,
16'h0DEB, 16'hFFFF,
16'h0DEC, 16'hFFFF,
16'h0DED, 16'hFFFF,
16'h0DEE, 16'hFFFF,
16'h0DEF, 16'hFFFF,
16'h0DF0, 16'hFFFF,
16'h0DF1, 16'hFFFF,
16'h0DF2, 16'hFFFF,
16'h0DF3, 16'hFFFF,
16'h0DF4, 16'hFFFF,
16'h0DF5, 16'hFFFF,
16'h0DF6, 16'hFFFF,
16'h0DF7, 16'hFFFF,
16'h0DF8, 16'hFFFF,
16'h0DF9, 16'hFFFF,
16'h0DFA, 16'hFFFF,
16'h0DFB, 16'hFFFF,
16'h0DFC, 16'hFFFF,
16'h0DFD, 16'hFFFF,
16'h0DFE, 16'hFFFF,
16'h0DFF, 16'hFFFF,
16'h0E00, 16'hFFFF,
16'h0E01, 16'hFFFF,
16'h0E02, 16'hFFFF,
16'h0E03, 16'hFFFF,
16'h0E04, 16'hFFFF,
16'h0E05, 16'hFFFF,
16'h0E06, 16'hFFFF,
16'h0E07, 16'hFFFF,
16'h0E08, 16'hFFFF,
16'h0E09, 16'hFFFF,
16'h0E0A, 16'hFFFF,
16'h0E0B, 16'hFFFF,
16'h0E0C, 16'hFFFF,
16'h0E0D, 16'hFFFF,
16'h0E0E, 16'hFFFF,
16'h0E0F, 16'hFFFF,
16'h0E10, 16'hFFFF,
16'h0E11, 16'hFFFF,
16'h0E12, 16'hFFFF,
16'h0E13, 16'hFFFF,
16'h0E14, 16'hFFFF,
16'h0E15, 16'hFFFF,
16'h0E16, 16'hFFFF,
16'h0E17, 16'hFFFF,
16'h0E18, 16'hFFFF,
16'h0E19, 16'hFFFF,
16'h0E1A, 16'hFFFF,
16'h0E1B, 16'hFFFF,
16'h0E1C, 16'hFFFF,
16'h0E1D, 16'hFFFF,
16'h0E1E, 16'hFFFF,
16'h0E1F, 16'hFFFF,
16'h0E20, 16'hFFFF,
16'h0E21, 16'hFFFF,
16'h0E22, 16'hFFFF,
16'h0E23, 16'hFFFF,
16'h0E24, 16'hFFFF,
16'h0E25, 16'hFFFF,
16'h0E26, 16'hFFFF,
16'h0E27, 16'hFFFF,
16'h0E28, 16'hFFFF,
16'h0E29, 16'hFFFF,
16'h0E2A, 16'hFFFF,
16'h0E2B, 16'hFFFF,
16'h0E2C, 16'hFFFF,
16'h0E2D, 16'hFFFF,
16'h0E2E, 16'hFFFF,
16'h0E2F, 16'hFFFF,
16'h0E30, 16'hFFFF,
16'h0E31, 16'hFFFF,
16'h0E32, 16'hFFFF,
16'h0E33, 16'hFFFF,
16'h0E34, 16'hFFFF,
16'h0E35, 16'hFFFF,
16'h0E36, 16'hFFFF,
16'h0E37, 16'hFFFF,
16'h0E38, 16'hFFFF,
16'h0E39, 16'hFFFF,
16'h0E3A, 16'hFFFF,
16'h0E3B, 16'hFFFF,
16'h0E3C, 16'hFFFF,
16'h0E3D, 16'hFFFF,
16'h0E3E, 16'hFFFF,
16'h0E3F, 16'hFFFF,
16'h0E40, 16'hFFFF,
16'h0E41, 16'hFFFF,
16'h0E42, 16'hFFFF,
16'h0E43, 16'hFFFF,
16'h0E44, 16'hFFFF,
16'h0E45, 16'hFFFF,
16'h0E46, 16'hFFFF,
16'h0E47, 16'hFFFF,
16'h0E48, 16'hFFFF,
16'h0E49, 16'hFFFF,
16'h0E4A, 16'hFFFF,
16'h0E4B, 16'hFFFF,
16'h0E4C, 16'hFFFF,
16'h0E4D, 16'hFFFF,
16'h0E4E, 16'hFFFF,
16'h0E4F, 16'hFFFF,
16'h0E50, 16'hFFFF,
16'h0E51, 16'hFFFF,
16'h0E52, 16'hFFFF,
16'h0E53, 16'hFFFF,
16'h0E54, 16'hFFFF,
16'h0E55, 16'hFFFF,
16'h0E56, 16'hFFFF,
16'h0E57, 16'hFFFF,
16'h0E58, 16'hFFFF,
16'h0E59, 16'hFFFF,
16'h0E5A, 16'hFFFF,
16'h0E5B, 16'hFFFF,
16'h0E5C, 16'hFFFF,
16'h0E5D, 16'hFFFF,
16'h0E5E, 16'hFFFF,
16'h0E5F, 16'hFFFF,
16'h0E60, 16'hFFFF,
16'h0E61, 16'hFFFF,
16'h0E62, 16'hFFFF,
16'h0E63, 16'hFFFF,
16'h0E64, 16'hFFFF,
16'h0E65, 16'hFFFF,
16'h0E66, 16'hFFFF,
16'h0E67, 16'hFFFF,
16'h0E68, 16'hFFFF,
16'h0E69, 16'hFFFF,
16'h0E6A, 16'hFFFF,
16'h0E6B, 16'hFFFF,
16'h0E6C, 16'hFFFF,
16'h0E6D, 16'hFFFF,
16'h0E6E, 16'hFFFF,
16'h0E6F, 16'hFFFF,
16'h0E70, 16'hFFFF,
16'h0E71, 16'hFFFF,
16'h0E72, 16'hFFFF,
16'h0E73, 16'hFFFF,
16'h0E74, 16'hFFFF,
16'h0E75, 16'hFFFF,
16'h0E76, 16'hFFFF,
16'h0E77, 16'hFFFF,
16'h0E78, 16'hFFFF,
16'h0E79, 16'hFFFF,
16'h0E7A, 16'hFFFF,
16'h0E7B, 16'hFFFF,
16'h0E7C, 16'hFFFF,
16'h0E7D, 16'hFFFF,
16'h0E7E, 16'hFFFF,
16'h0E7F, 16'hFFFF,
16'h0E80, 16'hFFFF,
16'h0E81, 16'hFFFF,
16'h0E82, 16'hFFFF,
16'h0E83, 16'hFFFF,
16'h0E84, 16'hFFFF,
16'h0E85, 16'hFFFF,
16'h0E86, 16'hFFFF,
16'h0E87, 16'hFFFF,
16'h0E88, 16'hFFFF,
16'h0E89, 16'hFFFF,
16'h0E8A, 16'hFFFF,
16'h0E8B, 16'hFFFF,
16'h0E8C, 16'hFFFF,
16'h0E8D, 16'hFFFF,
16'h0E8E, 16'hFFFF,
16'h0E8F, 16'hFFFF,
16'h0E90, 16'hFFFF,
16'h0E91, 16'hFFFF,
16'h0E92, 16'hFFFF,
16'h0E93, 16'hFFFF,
16'h0E94, 16'hFFFF,
16'h0E95, 16'hFFFF,
16'h0E96, 16'hFFFF,
16'h0E97, 16'hFFFF,
16'h0E98, 16'hFFFF,
16'h0E99, 16'hFFFF,
16'h0E9A, 16'hFFFF,
16'h0E9B, 16'hFFFF,
16'h0E9C, 16'hFFFF,
16'h0E9D, 16'hFFFF,
16'h0E9E, 16'hFFFF,
16'h0E9F, 16'hFFFF,
16'h0EA0, 16'hFFFF,
16'h0EA1, 16'hFFFF,
16'h0EA2, 16'hFFFF,
16'h0EA3, 16'hFFFF,
16'h0EA4, 16'hFFFF,
16'h0EA5, 16'hFFFF,
16'h0EA6, 16'hFFFF,
16'h0EA7, 16'hFFFF,
16'h0EA8, 16'hFFFF,
16'h0EA9, 16'hFFFF,
16'h0EAA, 16'hFFFF,
16'h0EAB, 16'hFFFF,
16'h0EAC, 16'hFFFF,
16'h0EAD, 16'hFFFF,
16'h0EAE, 16'hFFFF,
16'h0EAF, 16'hFFFF,
16'h0EB0, 16'hFFFF,
16'h0EB1, 16'hFFFF,
16'h0EB2, 16'hFFFF,
16'h0EB3, 16'hFFFF,
16'h0EB4, 16'hFFFF,
16'h0EB5, 16'hFFFF,
16'h0EB6, 16'hFFFF,
16'h0EB7, 16'hFFFF,
16'h0EB8, 16'hFFFF,
16'h0EB9, 16'hFFFF,
16'h0EBA, 16'hFFFF,
16'h0EBB, 16'hFFFF,
16'h0EBC, 16'hFFFF,
16'h0EBD, 16'hFFFF,
16'h0EBE, 16'hFFFF,
16'h0EBF, 16'hFFFF,
16'h0EC0, 16'hFFFF,
16'h0EC1, 16'hFFFF,
16'h0EC2, 16'hFFFF,
16'h0EC3, 16'hFFFF,
16'h0EC4, 16'hFFFF,
16'h0EC5, 16'hFFFF,
16'h0EC6, 16'hFFFF,
16'h0EC7, 16'hFFFF,
16'h0EC8, 16'hFFFF,
16'h0EC9, 16'hFFFF,
16'h0ECA, 16'hFFFF,
16'h0ECB, 16'hFFFF,
16'h0ECC, 16'hFFFF,
16'h0ECD, 16'hFFFF,
16'h0ECE, 16'hFFFF,
16'h0ECF, 16'hFFFF,
16'h0ED0, 16'hFFFF,
16'h0ED1, 16'hFFFF,
16'h0ED2, 16'hFFFF,
16'h0ED3, 16'hFFFF,
16'h0ED4, 16'hFFFF,
16'h0ED5, 16'hFFFF,
16'h0ED6, 16'hFFFF,
16'h0ED7, 16'hFFFF,
16'h0ED8, 16'hFFFF,
16'h0ED9, 16'hFFFF,
16'h0EDA, 16'hFFFF,
16'h0EDB, 16'hFFFF,
16'h0EDC, 16'hFFFF,
16'h0EDD, 16'hFFFF,
16'h0EDE, 16'hFFFF,
16'h0EDF, 16'hFFFF,
16'h0EE0, 16'hFFFF,
16'h0EE1, 16'hFFFF,
16'h0EE2, 16'hFFFF,
16'h0EE3, 16'hFFFF,
16'h0EE4, 16'hFFFF,
16'h0EE5, 16'hFFFF,
16'h0EE6, 16'hFFFF,
16'h0EE7, 16'hFFFF,
16'h0EE8, 16'hFFFF,
16'h0EE9, 16'hFFFF,
16'h0EEA, 16'hFFFF,
16'h0EEB, 16'hFFFF,
16'h0EEC, 16'hFFFF,
16'h0EED, 16'hFFFF,
16'h0EEE, 16'hFFFF,
16'h0EEF, 16'hFFFF,
16'h0EF0, 16'hFFFF,
16'h0EF1, 16'hFFFF,
16'h0EF2, 16'hFFFF,
16'h0EF3, 16'hFFFF,
16'h0EF4, 16'hFFFF,
16'h0EF5, 16'hFFFF,
16'h0EF6, 16'hFFFF,
16'h0EF7, 16'hFFFF,
16'h0EF8, 16'hFFFF,
16'h0EF9, 16'hFFFF,
16'h0EFA, 16'hFFFF,
16'h0EFB, 16'hFFFF,
16'h0EFC, 16'hFFFF,
16'h0EFD, 16'hFFFF,
16'h0EFE, 16'hFFFF,
16'h0EFF, 16'hFFFF,
16'h0F00, 16'hFFFF,
16'h0F01, 16'hFFFF,
16'h0F02, 16'hFFFF,
16'h0F03, 16'hFFFF,
16'h0F04, 16'hFFFF,
16'h0F05, 16'hFFFF,
16'h0F06, 16'hFFFF,
16'h0F07, 16'hFFFF,
16'h0F08, 16'hFFFF,
16'h0F09, 16'hFFFF,
16'h0F0A, 16'hFFFF,
16'h0F0B, 16'hFFFF,
16'h0F0C, 16'hFFFF,
16'h0F0D, 16'hFFFF,
16'h0F0E, 16'hFFFF,
16'h0F0F, 16'hFFFF,
16'h0F10, 16'hFFFF,
16'h0F11, 16'hFFFF,
16'h0F12, 16'hFFFF,
16'h0F13, 16'hFFFF,
16'h0F14, 16'hFFFF,
16'h0F15, 16'hFFFF,
16'h0F16, 16'hFFFF,
16'h0F17, 16'hFFFF,
16'h0F18, 16'hFFFF,
16'h0F19, 16'hFFFF,
16'h0F1A, 16'hFFFF,
16'h0F1B, 16'hFFFF,
16'h0F1C, 16'hFFFF,
16'h0F1D, 16'hFFFF,
16'h0F1E, 16'hFFFF,
16'h0F1F, 16'hFFFF,
16'h0F20, 16'hFFFF,
16'h0F21, 16'hFFFF,
16'h0F22, 16'hFFFF,
16'h0F23, 16'hFFFF,
16'h0F24, 16'hFFFF,
16'h0F25, 16'hFFFF,
16'h0F26, 16'hFFFF,
16'h0F27, 16'hFFFF,
16'h0F28, 16'hFFFF,
16'h0F29, 16'hFFFF,
16'h0F2A, 16'hFFFF,
16'h0F2B, 16'hFFFF,
16'h0F2C, 16'hFFFF,
16'h0F2D, 16'hFFFF,
16'h0F2E, 16'hFFFF,
16'h0F2F, 16'hFFFF,
16'h0F30, 16'hFFFF,
16'h0F31, 16'hFFFF,
16'h0F32, 16'hFFFF,
16'h0F33, 16'hFFFF,
16'h0F34, 16'hFFFF,
16'h0F35, 16'hFFFF,
16'h0F36, 16'hFFFF,
16'h0F37, 16'hFFFF,
16'h0F38, 16'hFFFF,
16'h0F39, 16'hFFFF,
16'h0F3A, 16'hFFFF,
16'h0F3B, 16'hFFFF,
16'h0F3C, 16'hFFFF,
16'h0F3D, 16'hFFFF,
16'h0F3E, 16'hFFFF,
16'h0F3F, 16'hFFFF,
16'h0F40, 16'hFFFF,
16'h0F41, 16'hFFFF,
16'h0F42, 16'hFFFF,
16'h0F43, 16'hFFFF,
16'h0F44, 16'hFFFF,
16'h0F45, 16'hFFFF,
16'h0F46, 16'hFFFF,
16'h0F47, 16'hFFFF,
16'h0F48, 16'hFFFF,
16'h0F49, 16'hFFFF,
16'h0F4A, 16'hFFFF,
16'h0F4B, 16'hFFFF,
16'h0F4C, 16'hFFFF,
16'h0F4D, 16'hFFFF,
16'h0F4E, 16'hFFFF,
16'h0F4F, 16'hFFFF,
16'h0F50, 16'hFFFF,
16'h0F51, 16'hFFFF,
16'h0F52, 16'hFFFF,
16'h0F53, 16'hFFFF,
16'h0F54, 16'hFFFF,
16'h0F55, 16'hFFFF,
16'h0F56, 16'hFFFF,
16'h0F57, 16'hFFFF,
16'h0F58, 16'hFFFF,
16'h0F59, 16'hFFFF,
16'h0F5A, 16'hFFFF,
16'h0F5B, 16'hFFFF,
16'h0F5C, 16'hFFFF,
16'h0F5D, 16'hFFFF,
16'h0F5E, 16'hFFFF,
16'h0F5F, 16'hFFFF,
16'h0F60, 16'hFFFF,
16'h0F61, 16'hFFFF,
16'h0F62, 16'hFFFF,
16'h0F63, 16'hFFFF,
16'h0F64, 16'hFFFF,
16'h0F65, 16'hFFFF,
16'h0F66, 16'hFFFF,
16'h0F67, 16'hFFFF,
16'h0F68, 16'hFFFF,
16'h0F69, 16'hFFFF,
16'h0F6A, 16'hFFFF,
16'h0F6B, 16'hFFFF,
16'h0F6C, 16'hFFFF,
16'h0F6D, 16'hFFFF,
16'h0F6E, 16'hFFFF,
16'h0F6F, 16'hFFFF,
16'h0F70, 16'hFFFF,
16'h0F71, 16'hFFFF,
16'h0F72, 16'hFFFF,
16'h0F73, 16'hFFFF,
16'h0F74, 16'hFFFF,
16'h0F75, 16'hFFFF,
16'h0F76, 16'hFFFF,
16'h0F77, 16'hFFFF,
16'h0F78, 16'hFFFF,
16'h0F79, 16'hFFFF,
16'h0F7A, 16'hFFFF,
16'h0F7B, 16'hFFFF,
16'h0F7C, 16'hFFFF,
16'h0F7D, 16'hFFFF,
16'h0F7E, 16'hFFFF,
16'h0F7F, 16'hFFFF,
16'h0F80, 16'hFFFF,
16'h0F81, 16'hFFFF,
16'h0F82, 16'hFFFF,
16'h0F83, 16'hFFFF,
16'h0F84, 16'hFFFF,
16'h0F85, 16'hFFFF,
16'h0F86, 16'hFFFF,
16'h0F87, 16'hFFFF,
16'h0F88, 16'hFFFF,
16'h0F89, 16'hFFFF,
16'h0F8A, 16'hFFFF,
16'h0F8B, 16'hFFFF,
16'h0F8C, 16'hFFFF,
16'h0F8D, 16'hFFFF,
16'h0F8E, 16'hFFFF,
16'h0F8F, 16'hFFFF,
16'h0F90, 16'hFFFF,
16'h0F91, 16'hFFFF,
16'h0F92, 16'hFFFF,
16'h0F93, 16'hFFFF,
16'h0F94, 16'hFFFF,
16'h0F95, 16'hFFFF,
16'h0F96, 16'hFFFF,
16'h0F97, 16'hFFFF,
16'h0F98, 16'hFFFF,
16'h0F99, 16'hFFFF,
16'h0F9A, 16'hFFFF,
16'h0F9B, 16'hFFFF,
16'h0F9C, 16'hFFFF,
16'h0F9D, 16'hFFFF,
16'h0F9E, 16'hFFFF,
16'h0F9F, 16'hFFFF,
16'h0FA0, 16'hFFFF,
16'h0FA1, 16'hFFFF,
16'h0FA2, 16'hFFFF,
16'h0FA3, 16'hFFFF,
16'h0FA4, 16'hFFFF,
16'h0FA5, 16'hFFFF,
16'h0FA6, 16'hFFFF,
16'h0FA7, 16'hFFFF,
16'h0FA8, 16'hFFFF,
16'h0FA9, 16'hFFFF,
16'h0FAA, 16'hFFFF,
16'h0FAB, 16'hFFFF,
16'h0FAC, 16'hFFFF,
16'h0FAD, 16'hFFFF,
16'h0FAE, 16'hFFFF,
16'h0FAF, 16'hFFFF,
16'h0FB0, 16'hFFFF,
16'h0FB1, 16'hFFFF,
16'h0FB2, 16'hFFFF,
16'h0FB3, 16'hFFFF,
16'h0FB4, 16'hFFFF,
16'h0FB5, 16'hFFFF,
16'h0FB6, 16'hFFFF,
16'h0FB7, 16'hFFFF,
16'h0FB8, 16'hFFFF,
16'h0FB9, 16'hFFFF,
16'h0FBA, 16'hFFFF,
16'h0FBB, 16'hFFFF,
16'h0FBC, 16'hFFFF,
16'h0FBD, 16'hFFFF,
16'h0FBE, 16'hFFFF,
16'h0FBF, 16'hFFFF,
16'h0FC0, 16'hFFFF,
16'h0FC1, 16'hFFFF,
16'h0FC2, 16'hFFFF,
16'h0FC3, 16'hFFFF,
16'h0FC4, 16'hFFFF,
16'h0FC5, 16'hFFFF,
16'h0FC6, 16'hFFFF,
16'h0FC7, 16'hFFFF,
16'h0FC8, 16'hFFFF,
16'h0FC9, 16'hFFFF,
16'h0FCA, 16'hFFFF,
16'h0FCB, 16'hFFFF,
16'h0FCC, 16'hFFFF,
16'h0FCD, 16'hFFFF,
16'h0FCE, 16'hFFFF,
16'h0FCF, 16'hFFFF,
16'h0FD0, 16'hFFFF,
16'h0FD1, 16'hFFFF,
16'h0FD2, 16'hFFFF,
16'h0FD3, 16'hFFFF,
16'h0FD4, 16'hFFFF,
16'h0FD5, 16'hFFFF,
16'h0FD6, 16'hFFFF,
16'h0FD7, 16'hFFFF,
16'h0FD8, 16'hFFFF,
16'h0FD9, 16'hFFFF,
16'h0FDA, 16'hFFFF,
16'h0FDB, 16'hFFFF,
16'h0FDC, 16'hFFFF,
16'h0FDD, 16'hFFFF,
16'h0FDE, 16'hFFFF,
16'h0FDF, 16'hFFFF,
16'h0FE0, 16'hFFFF,
16'h0FE1, 16'hFFFF,
16'h0FE2, 16'hFFFF,
16'h0FE3, 16'hFFFF,
16'h0FE4, 16'hFFFF,
16'h0FE5, 16'hFFFF,
16'h0FE6, 16'hFFFF,
16'h0FE7, 16'hFFFF,
16'h0FE8, 16'hFFFF,
16'h0FE9, 16'hFFFF,
16'h0FEA, 16'hFFFF,
16'h0FEB, 16'hFFFF,
16'h0FEC, 16'hFFFF,
16'h0FED, 16'hFFFF,
16'h0FEE, 16'hFFFF,
16'h0FEF, 16'hFFFF,
16'h0FF0, 16'hFFFF,
16'h0FF1, 16'hFFFF,
16'h0FF2, 16'hFFFF,
16'h0FF3, 16'hFFFF,
16'h0FF4, 16'hFFFF,
16'h0FF5, 16'hFFFF,
16'h0FF6, 16'hFFFF,
16'h0FF7, 16'hFFFF,
16'h0FF8, 16'hFFFF,
16'h0FF9, 16'hFFFF,
16'h0FFA, 16'hFFFF,
16'h0FFB, 16'hFFFF,
16'h0FFC, 16'hFFFF,
16'h0FFD, 16'hFFFF,
16'h0FFE, 16'hFFFF,
16'h0FFF, 16'hFFFF,
16'h1000, 16'hFFFF,
16'h1001, 16'hFFFF,
16'h1002, 16'hFFFF,
16'h1003, 16'hFFFF,
16'h1004, 16'hFFFF,
16'h1005, 16'hFFFF,
16'h1006, 16'hFFFF,
16'h1007, 16'hFFFF,
16'h1008, 16'hFFFF,
16'h1009, 16'hFFFF,
16'h100A, 16'hFFFF,
16'h100B, 16'hFFFF,
16'h100C, 16'hFFFF,
16'h100D, 16'hFFFF,
16'h100E, 16'hFFFF,
16'h100F, 16'hFFFF,
16'h1010, 16'hFFFF,
16'h1011, 16'hFFFF,
16'h1012, 16'hFFFF,
16'h1013, 16'hFFFF,
16'h1014, 16'hFFFF,
16'h1015, 16'hFFFF,
16'h1016, 16'hFFFF,
16'h1017, 16'hFFFF,
16'h1018, 16'hFFFF,
16'h1019, 16'hFFFF,
16'h101A, 16'hFFFF,
16'h101B, 16'hFFFF,
16'h101C, 16'hFFFF,
16'h101D, 16'hFFFF,
16'h101E, 16'hFFFF,
16'h101F, 16'hFFFF,
16'h1020, 16'hFFFF,
16'h1021, 16'hFFFF,
16'h1022, 16'hFFFF,
16'h1023, 16'hFFFF,
16'h1024, 16'hFFFF,
16'h1025, 16'hFFFF,
16'h1026, 16'hFFFF,
16'h1027, 16'hFFFF,
16'h1028, 16'hFFFF,
16'h1029, 16'hFFFF,
16'h102A, 16'hFFFF,
16'h102B, 16'hFFFF,
16'h102C, 16'hFFFF,
16'h102D, 16'hFFFF,
16'h102E, 16'hFFFF,
16'h102F, 16'hFFFF,
16'h1030, 16'hFFFF,
16'h1031, 16'hFFFF,
16'h1032, 16'hFFFF,
16'h1033, 16'hFFFF,
16'h1034, 16'hFFFF,
16'h1035, 16'hFFFF,
16'h1036, 16'hFFFF,
16'h1037, 16'hFFFF,
16'h1038, 16'hFFFF,
16'h1039, 16'hFFFF,
16'h103A, 16'hFFFF,
16'h103B, 16'hFFFF,
16'h103C, 16'hFFFF,
16'h103D, 16'hFFFF,
16'h103E, 16'hFFFF,
16'h103F, 16'hFFFF,
16'h1040, 16'hFFFF,
16'h1041, 16'hFFFF,
16'h1042, 16'hFFFF,
16'h1043, 16'hFFFF,
16'h1044, 16'hFFFF,
16'h1045, 16'hFFFF,
16'h1046, 16'hFFFF,
16'h1047, 16'hFFFF,
16'h1048, 16'hFFFF,
16'h1049, 16'hFFFF,
16'h104A, 16'hFFFF,
16'h104B, 16'hFFFF,
16'h104C, 16'hFFFF,
16'h104D, 16'hFFFF,
16'h104E, 16'hFFFF,
16'h104F, 16'hFFFF,
16'h1050, 16'hFFFF,
16'h1051, 16'hFFFF,
16'h1052, 16'hFFFF,
16'h1053, 16'hFFFF,
16'h1054, 16'hFFFF,
16'h1055, 16'hFFFF,
16'h1056, 16'hFFFF,
16'h1057, 16'hFFFF,
16'h1058, 16'hFFFF,
16'h1059, 16'hFFFF,
16'h105A, 16'hFFFF,
16'h105B, 16'hFFFF,
16'h105C, 16'hFFFF,
16'h105D, 16'hFFFF,
16'h105E, 16'hFFFF,
16'h105F, 16'hFFFF,
16'h1060, 16'hFFFF,
16'h1061, 16'hFFFF,
16'h1062, 16'hFFFF,
16'h1063, 16'hFFFF,
16'h1064, 16'hFFFF,
16'h1065, 16'hFFFF,
16'h1066, 16'hFFFF,
16'h1067, 16'hFFFF,
16'h1068, 16'hFFFF,
16'h1069, 16'hFFFF,
16'h106A, 16'hFFFF,
16'h106B, 16'hFFFF,
16'h106C, 16'hFFFF,
16'h106D, 16'hFFFF,
16'h106E, 16'hFFFF,
16'h106F, 16'hFFFF,
16'h1070, 16'hFFFF,
16'h1071, 16'hFFFF,
16'h1072, 16'hFFFF,
16'h1073, 16'hFFFF,
16'h1074, 16'hFFFF,
16'h1075, 16'hFFFF,
16'h1076, 16'hFFFF,
16'h1077, 16'hFFFF,
16'h1078, 16'hFFFF,
16'h1079, 16'hFFFF,
16'h107A, 16'hFFFF,
16'h107B, 16'hFFFF,
16'h107C, 16'hFFFF,
16'h107D, 16'hFFFF,
16'h107E, 16'hFFFF,
16'h107F, 16'hFFFF,
16'h1080, 16'hFFFF,
16'h1081, 16'hFFFF,
16'h1082, 16'hFFFF,
16'h1083, 16'hFFFF,
16'h1084, 16'hFFFF,
16'h1085, 16'hFFFF,
16'h1086, 16'hFFFF,
16'h1087, 16'hFFFF,
16'h1088, 16'hFFFF,
16'h1089, 16'hFFFF,
16'h108A, 16'hFFFF,
16'h108B, 16'hFFFF,
16'h108C, 16'hFFFF,
16'h108D, 16'hFFFF,
16'h108E, 16'hFFFF,
16'h108F, 16'hFFFF,
16'h1090, 16'hFFFF,
16'h1091, 16'hFFFF,
16'h1092, 16'hFFFF,
16'h1093, 16'hFFFF,
16'h1094, 16'hFFFF,
16'h1095, 16'hFFFF,
16'h1096, 16'hFFFF,
16'h1097, 16'hFFFF,
16'h1098, 16'hFFFF,
16'h1099, 16'hFFFF,
16'h109A, 16'hFFFF,
16'h109B, 16'hFFFF,
16'h109C, 16'hFFFF,
16'h109D, 16'hFFFF,
16'h109E, 16'hFFFF,
16'h109F, 16'hFFFF,
16'h10A0, 16'hFFFF,
16'h10A1, 16'hFFFF,
16'h10A2, 16'hFFFF,
16'h10A3, 16'hFFFF,
16'h10A4, 16'hFFFF,
16'h10A5, 16'hFFFF,
16'h10A6, 16'hFFFF,
16'h10A7, 16'hFFFF,
16'h10A8, 16'hFFFF,
16'h10A9, 16'hFFFF,
16'h10AA, 16'hFFFF,
16'h10AB, 16'hFFFF,
16'h10AC, 16'hFFFF,
16'h10AD, 16'hFFFF,
16'h10AE, 16'hFFFF,
16'h10AF, 16'hFFFF,
16'h10B0, 16'hFFFF,
16'h10B1, 16'hFFFF,
16'h10B2, 16'hFFFF,
16'h10B3, 16'hFFFF,
16'h10B4, 16'hFFFF,
16'h10B5, 16'hFFFF,
16'h10B6, 16'hFFFF,
16'h10B7, 16'hFFFF,
16'h10B8, 16'hFFFF,
16'h10B9, 16'hFFFF,
16'h10BA, 16'hFFFF,
16'h10BB, 16'hFFFF,
16'h10BC, 16'hFFFF,
16'h10BD, 16'hFFFF,
16'h10BE, 16'hFFFF,
16'h10BF, 16'hFFFF,
16'h10C0, 16'hFFFF,
16'h10C1, 16'hFFFF,
16'h10C2, 16'hFFFF,
16'h10C3, 16'hFFFF,
16'h10C4, 16'hFFFF,
16'h10C5, 16'hFFFF,
16'h10C6, 16'hFFFF,
16'h10C7, 16'hFFFF,
16'h10C8, 16'hFFFF,
16'h10C9, 16'hFFFF,
16'h10CA, 16'hFFFF,
16'h10CB, 16'hFFFF,
16'h10CC, 16'hFFFF,
16'h10CD, 16'hFFFF,
16'h10CE, 16'hFFFF,
16'h10CF, 16'hFFFF,
16'h10D0, 16'hFFFF,
16'h10D1, 16'hFFFF,
16'h10D2, 16'hFFFF,
16'h10D3, 16'hFFFF,
16'h10D4, 16'hFFFF,
16'h10D5, 16'hFFFF,
16'h10D6, 16'hFFFF,
16'h10D7, 16'hFFFF,
16'h10D8, 16'hFFFF,
16'h10D9, 16'hFFFF,
16'h10DA, 16'hFFFF,
16'h10DB, 16'hFFFF,
16'h10DC, 16'hFFFF,
16'h10DD, 16'hFFFF,
16'h10DE, 16'hFFFF,
16'h10DF, 16'hFFFF,
16'h10E0, 16'hFFFF,
16'h10E1, 16'hFFFF,
16'h10E2, 16'hFFFF,
16'h10E3, 16'hFFFF,
16'h10E4, 16'hFFFF,
16'h10E5, 16'hFFFF,
16'h10E6, 16'hFFFF,
16'h10E7, 16'hFFFF,
16'h10E8, 16'hFFFF,
16'h10E9, 16'hFFFF,
16'h10EA, 16'hFFFF,
16'h10EB, 16'hFFFF,
16'h10EC, 16'hFFFF,
16'h10ED, 16'hFFFF,
16'h10EE, 16'hFFFF,
16'h10EF, 16'hFFFF,
16'h10F0, 16'hFFFF,
16'h10F1, 16'hFFFF,
16'h10F2, 16'hFFFF,
16'h10F3, 16'hFFFF,
16'h10F4, 16'hFFFF,
16'h10F5, 16'hFFFF,
16'h10F6, 16'hFFFF,
16'h10F7, 16'hFFFF,
16'h10F8, 16'hFFFF,
16'h10F9, 16'hFFFF,
16'h10FA, 16'hFFFF,
16'h10FB, 16'hFFFF,
16'h10FC, 16'hFFFF,
16'h10FD, 16'hFFFF,
16'h10FE, 16'hFFFF,
16'h10FF, 16'hFFFF,
16'h1100, 16'hFFFF,
16'h1101, 16'hFFFF,
16'h1102, 16'hFFFF,
16'h1103, 16'hFFFF,
16'h1104, 16'hFFFF,
16'h1105, 16'hFFFF,
16'h1106, 16'hFFFF,
16'h1107, 16'hFFFF,
16'h1108, 16'hFFFF,
16'h1109, 16'hFFFF,
16'h110A, 16'hFFFF,
16'h110B, 16'hFFFF,
16'h110C, 16'hFFFF,
16'h110D, 16'hFFFF,
16'h110E, 16'hFFFF,
16'h110F, 16'hFFFF,
16'h1110, 16'hFFFF,
16'h1111, 16'hFFFF,
16'h1112, 16'hFFFF,
16'h1113, 16'hFFFF,
16'h1114, 16'hFFFF,
16'h1115, 16'hFFFF,
16'h1116, 16'hFFFF,
16'h1117, 16'hFFFF,
16'h1118, 16'hFFFF,
16'h1119, 16'hFFFF,
16'h111A, 16'hFFFF,
16'h111B, 16'hFFFF,
16'h111C, 16'hFFFF,
16'h111D, 16'hFFFF,
16'h111E, 16'hFFFF,
16'h111F, 16'hFFFF,
16'h1120, 16'hFFFF,
16'h1121, 16'hFFFF,
16'h1122, 16'hFFFF,
16'h1123, 16'hFFFF,
16'h1124, 16'hFFFF,
16'h1125, 16'hFFFF,
16'h1126, 16'hFFFF,
16'h1127, 16'hFFFF,
16'h1128, 16'hFFFF,
16'h1129, 16'hFFFF,
16'h112A, 16'hFFFF,
16'h112B, 16'hFFFF,
16'h112C, 16'hFFFF,
16'h112D, 16'hFFFF,
16'h112E, 16'hFFFF,
16'h112F, 16'hFFFF,
16'h1130, 16'hFFFF,
16'h1131, 16'hFFFF,
16'h1132, 16'hFFFF,
16'h1133, 16'hFFFF,
16'h1134, 16'hFFFF,
16'h1135, 16'hFFFF,
16'h1136, 16'hFFFF,
16'h1137, 16'hFFFF,
16'h1138, 16'hFFFF,
16'h1139, 16'hFFFF,
16'h113A, 16'hFFFF,
16'h113B, 16'hFFFF,
16'h113C, 16'hFFFF,
16'h113D, 16'hFFFF,
16'h113E, 16'hFFFF,
16'h113F, 16'hFFFF,
16'h1140, 16'hFFFF,
16'h1141, 16'hFFFF,
16'h1142, 16'hFFFF,
16'h1143, 16'hFFFF,
16'h1144, 16'hFFFF,
16'h1145, 16'hFFFF,
16'h1146, 16'hFFFF,
16'h1147, 16'hFFFF,
16'h1148, 16'hFFFF,
16'h1149, 16'hFFFF,
16'h114A, 16'hFFFF,
16'h114B, 16'hFFFF,
16'h114C, 16'hFFFF,
16'h114D, 16'hFFFF,
16'h114E, 16'hFFFF,
16'h114F, 16'hFFFF,
16'h1150, 16'hFFFF,
16'h1151, 16'hFFFF,
16'h1152, 16'hFFFF,
16'h1153, 16'hFFFF,
16'h1154, 16'hFFFF,
16'h1155, 16'hFFFF,
16'h1156, 16'hFFFF,
16'h1157, 16'hFFFF,
16'h1158, 16'hFFFF,
16'h1159, 16'hFFFF,
16'h115A, 16'hFFFF,
16'h115B, 16'hFFFF,
16'h115C, 16'hFFFF,
16'h115D, 16'hFFFF,
16'h115E, 16'hFFFF,
16'h115F, 16'hFFFF,
16'h1160, 16'hFFFF,
16'h1161, 16'hFFFF,
16'h1162, 16'hFFFF,
16'h1163, 16'hFFFF,
16'h1164, 16'hFFFF,
16'h1165, 16'hFFFF,
16'h1166, 16'hFFFF,
16'h1167, 16'hFFFF,
16'h1168, 16'hFFFF,
16'h1169, 16'hFFFF,
16'h116A, 16'hFFFF,
16'h116B, 16'hFFFF,
16'h116C, 16'hFFFF,
16'h116D, 16'hFFFF,
16'h116E, 16'hFFFF,
16'h116F, 16'hFFFF,
16'h1170, 16'hFFFF,
16'h1171, 16'hFFFF,
16'h1172, 16'hFFFF,
16'h1173, 16'hFFFF,
16'h1174, 16'hFFFF,
16'h1175, 16'hFFFF,
16'h1176, 16'hFFFF,
16'h1177, 16'hFFFF,
16'h1178, 16'hFFFF,
16'h1179, 16'hFFFF,
16'h117A, 16'hFFFF,
16'h117B, 16'hFFFF,
16'h117C, 16'hFFFF,
16'h117D, 16'hFFFF,
16'h117E, 16'hFFFF,
16'h117F, 16'hFFFF,
16'h1180, 16'hFFFF,
16'h1181, 16'hFFFF,
16'h1182, 16'hFFFF,
16'h1183, 16'hFFFF,
16'h1184, 16'hFFFF,
16'h1185, 16'hFFFF,
16'h1186, 16'hFFFF,
16'h1187, 16'hFFFF,
16'h1188, 16'hFFFF,
16'h1189, 16'hFFFF,
16'h118A, 16'hFFFF,
16'h118B, 16'hFFFF,
16'h118C, 16'hFFFF,
16'h118D, 16'hFFFF,
16'h118E, 16'hFFFF,
16'h118F, 16'hFFFF,
16'h1190, 16'hFFFF,
16'h1191, 16'hFFFF,
16'h1192, 16'hFFFF,
16'h1193, 16'hFFFF,
16'h1194, 16'hFFFF,
16'h1195, 16'hFFFF,
16'h1196, 16'hFFFF,
16'h1197, 16'hFFFF,
16'h1198, 16'hFFFF,
16'h1199, 16'hFFFF,
16'h119A, 16'hFFFF,
16'h119B, 16'hFFFF,
16'h119C, 16'hFFFF,
16'h119D, 16'hFFFF,
16'h119E, 16'hFFFF,
16'h119F, 16'hFFFF,
16'h11A0, 16'hFFFF,
16'h11A1, 16'hFFFF,
16'h11A2, 16'hFFFF,
16'h11A3, 16'hFFFF,
16'h11A4, 16'hFFFF,
16'h11A5, 16'hFFFF,
16'h11A6, 16'hFFFF,
16'h11A7, 16'hFFFF,
16'h11A8, 16'hFFFF,
16'h11A9, 16'hFFFF,
16'h11AA, 16'hFFFF,
16'h11AB, 16'hFFFF,
16'h11AC, 16'hFFFF,
16'h11AD, 16'hFFFF,
16'h11AE, 16'hFFFF,
16'h11AF, 16'hFFFF,
16'h11B0, 16'hFFFF,
16'h11B1, 16'hFFFF,
16'h11B2, 16'hFFFF,
16'h11B3, 16'hFFFF,
16'h11B4, 16'hFFFF,
16'h11B5, 16'hFFFF,
16'h11B6, 16'hFFFF,
16'h11B7, 16'hFFFF,
16'h11B8, 16'hFFFF,
16'h11B9, 16'hFFFF,
16'h11BA, 16'hFFFF,
16'h11BB, 16'hFFFF,
16'h11BC, 16'hFFFF,
16'h11BD, 16'hFFFF,
16'h11BE, 16'hFFFF,
16'h11BF, 16'hFFFF,
16'h11C0, 16'hFFFF,
16'h11C1, 16'hFFFF,
16'h11C2, 16'hFFFF,
16'h11C3, 16'hFFFF,
16'h11C4, 16'hFFFF,
16'h11C5, 16'hFFFF,
16'h11C6, 16'hFFFF,
16'h11C7, 16'hFFFF,
16'h11C8, 16'hFFFF,
16'h11C9, 16'hFFFF,
16'h11CA, 16'hFFFF,
16'h11CB, 16'hFFFF,
16'h11CC, 16'hFFFF,
16'h11CD, 16'hFFFF,
16'h11CE, 16'hFFFF,
16'h11CF, 16'hFFFF,
16'h11D0, 16'hFFFF,
16'h11D1, 16'hFFFF,
16'h11D2, 16'hFFFF,
16'h11D3, 16'hFFFF,
16'h11D4, 16'hFFFF,
16'h11D5, 16'hFFFF,
16'h11D6, 16'hFFFF,
16'h11D7, 16'hFFFF,
16'h11D8, 16'hFFFF,
16'h11D9, 16'hFFFF,
16'h11DA, 16'hFFFF,
16'h11DB, 16'hFFFF,
16'h11DC, 16'hFFFF,
16'h11DD, 16'hFFFF,
16'h11DE, 16'hFFFF,
16'h11DF, 16'hFFFF,
16'h11E0, 16'hFFFF,
16'h11E1, 16'hFFFF,
16'h11E2, 16'hFFFF,
16'h11E3, 16'hFFFF,
16'h11E4, 16'hFFFF,
16'h11E5, 16'hFFFF,
16'h11E6, 16'hFFFF,
16'h11E7, 16'hFFFF,
16'h11E8, 16'hFFFF,
16'h11E9, 16'hFFFF,
16'h11EA, 16'hFFFF,
16'h11EB, 16'hFFFF,
16'h11EC, 16'hFFFF,
16'h11ED, 16'hFFFF,
16'h11EE, 16'hFFFF,
16'h11EF, 16'hFFFF,
16'h11F0, 16'hFFFF,
16'h11F1, 16'hFFFF,
16'h11F2, 16'hFFFF,
16'h11F3, 16'hFFFF,
16'h11F4, 16'hFFFF,
16'h11F5, 16'hFFFF,
16'h11F6, 16'hFFFF,
16'h11F7, 16'hFFFF,
16'h11F8, 16'hFFFF,
16'h11F9, 16'hFFFF,
16'h11FA, 16'hFFFF,
16'h11FB, 16'hFFFF,
16'h11FC, 16'hFFFF,
16'h11FD, 16'hFFFF,
16'h11FE, 16'hFFFF,
16'h11FF, 16'hFFFF,
16'h1200, 16'hFFFF,
16'h1201, 16'hFFFF,
16'h1202, 16'hFFFF,
16'h1203, 16'hFFFF,
16'h1204, 16'hFFFF,
16'h1205, 16'hFFFF,
16'h1206, 16'hFFFF,
16'h1207, 16'hFFFF,
16'h1208, 16'hFFFF,
16'h1209, 16'hFFFF,
16'h120A, 16'hFFFF,
16'h120B, 16'hFFFF,
16'h120C, 16'hFFFF,
16'h120D, 16'hFFFF,
16'h120E, 16'hFFFF,
16'h120F, 16'hFFFF,
16'h1210, 16'hFFFF,
16'h1211, 16'hFFFF,
16'h1212, 16'hFFFF,
16'h1213, 16'hFFFF,
16'h1214, 16'hFFFF,
16'h1215, 16'hFFFF,
16'h1216, 16'hFFFF,
16'h1217, 16'hFFFF,
16'h1218, 16'hFFFF,
16'h1219, 16'hFFFF,
16'h121A, 16'hFFFF,
16'h121B, 16'hFFFF,
16'h121C, 16'hFFFF,
16'h121D, 16'hFFFF,
16'h121E, 16'hFFFF,
16'h121F, 16'hFFFF,
16'h1220, 16'hFFFF,
16'h1221, 16'hFFFF,
16'h1222, 16'hFFFF,
16'h1223, 16'hFFFF,
16'h1224, 16'hFFFF,
16'h1225, 16'hFFFF,
16'h1226, 16'hFFFF,
16'h1227, 16'hFFFF,
16'h1228, 16'hFFFF,
16'h1229, 16'hFFFF,
16'h122A, 16'hFFFF,
16'h122B, 16'hFFFF,
16'h122C, 16'hFFFF,
16'h122D, 16'hFFFF,
16'h122E, 16'hFFFF,
16'h122F, 16'hFFFF,
16'h1230, 16'hFFFF,
16'h1231, 16'hFFFF,
16'h1232, 16'hFFFF,
16'h1233, 16'hFFFF,
16'h1234, 16'hFFFF,
16'h1235, 16'hFFFF,
16'h1236, 16'hFFFF,
16'h1237, 16'hFFFF,
16'h1238, 16'hFFFF,
16'h1239, 16'hFFFF,
16'h123A, 16'hFFFF,
16'h123B, 16'hFFFF,
16'h123C, 16'hFFFF,
16'h123D, 16'hFFFF,
16'h123E, 16'hFFFF,
16'h123F, 16'hFFFF,
16'h1240, 16'hFFFF,
16'h1241, 16'hFFFF,
16'h1242, 16'hFFFF,
16'h1243, 16'hFFFF,
16'h1244, 16'hFFFF,
16'h1245, 16'hFFFF,
16'h1246, 16'hFFFF,
16'h1247, 16'hFFFF,
16'h1248, 16'hFFFF,
16'h1249, 16'hFFFF,
16'h124A, 16'hFFFF,
16'h124B, 16'hFFFF,
16'h124C, 16'hFFFF,
16'h124D, 16'hFFFF,
16'h124E, 16'hFFFF,
16'h124F, 16'hFFFF,
16'h1250, 16'hFFFF,
16'h1251, 16'hFFFF,
16'h1252, 16'hFFFF,
16'h1253, 16'hFFFF,
16'h1254, 16'hFFFF,
16'h1255, 16'hFFFF,
16'h1256, 16'hFFFF,
16'h1257, 16'hFFFF,
16'h1258, 16'hFFFF,
16'h1259, 16'hFFFF,
16'h125A, 16'hFFFF,
16'h125B, 16'hFFFF,
16'h125C, 16'hFFFF,
16'h125D, 16'hFFFF,
16'h125E, 16'hFFFF,
16'h125F, 16'hFFFF,
16'h1260, 16'hFFFF,
16'h1261, 16'hFFFF,
16'h1262, 16'hFFFF,
16'h1263, 16'hFFFF,
16'h1264, 16'hFFFF,
16'h1265, 16'hFFFF,
16'h1266, 16'hFFFF,
16'h1267, 16'hFFFF,
16'h1268, 16'hFFFF,
16'h1269, 16'hFFFF,
16'h126A, 16'hFFFF,
16'h126B, 16'hFFFF,
16'h126C, 16'hFFFF,
16'h126D, 16'hFFFF,
16'h126E, 16'hFFFF,
16'h126F, 16'hFFFF,
16'h1270, 16'hFFFF,
16'h1271, 16'hFFFF,
16'h1272, 16'hFFFF,
16'h1273, 16'hFFFF,
16'h1274, 16'hFFFF,
16'h1275, 16'hFFFF,
16'h1276, 16'hFFFF,
16'h1277, 16'hFFFF,
16'h1278, 16'hFFFF,
16'h1279, 16'hFFFF,
16'h127A, 16'hFFFF,
16'h127B, 16'hFFFF,
16'h127C, 16'hFFFF,
16'h127D, 16'hFFFF,
16'h127E, 16'hFFFF,
16'h127F, 16'hFFFF,
16'h1280, 16'hFFFF,
16'h1281, 16'hFFFF,
16'h1282, 16'hFFFF,
16'h1283, 16'hFFFF,
16'h1284, 16'hFFFF,
16'h1285, 16'hFFFF,
16'h1286, 16'hFFFF,
16'h1287, 16'hFFFF,
16'h1288, 16'hFFFF,
16'h1289, 16'hFFFF,
16'h128A, 16'hFFFF,
16'h128B, 16'hFFFF,
16'h128C, 16'hFFFF,
16'h128D, 16'hFFFF,
16'h128E, 16'hFFFF,
16'h128F, 16'hFFFF,
16'h1290, 16'hFFFF,
16'h1291, 16'hFFFF,
16'h1292, 16'hFFFF,
16'h1293, 16'hFFFF,
16'h1294, 16'hFFFF,
16'h1295, 16'hFFFF,
16'h1296, 16'hFFFF,
16'h1297, 16'hFFFF,
16'h1298, 16'hFFFF,
16'h1299, 16'hFFFF,
16'h129A, 16'hFFFF,
16'h129B, 16'hFFFF,
16'h129C, 16'hFFFF,
16'h129D, 16'hFFFF,
16'h129E, 16'hFFFF,
16'h129F, 16'hFFFF,
16'h12A0, 16'hFFFF,
16'h12A1, 16'hFFFF,
16'h12A2, 16'hFFFF,
16'h12A3, 16'hFFFF,
16'h12A4, 16'hFFFF,
16'h12A5, 16'hFFFF,
16'h12A6, 16'hFFFF,
16'h12A7, 16'hFFFF,
16'h12A8, 16'hFFFF,
16'h12A9, 16'hFFFF,
16'h12AA, 16'hFFFF,
16'h12AB, 16'hFFFF,
16'h12AC, 16'hFFFF,
16'h12AD, 16'hFFFF,
16'h12AE, 16'hFFFF,
16'h12AF, 16'hFFFF,
16'h12B0, 16'hFFFF,
16'h12B1, 16'hFFFF,
16'h12B2, 16'hFFFF,
16'h12B3, 16'hFFFF,
16'h12B4, 16'hFFFF,
16'h12B5, 16'hFFFF,
16'h12B6, 16'hFFFF,
16'h12B7, 16'hFFFF,
16'h12B8, 16'hFFFF,
16'h12B9, 16'hFFFF,
16'h12BA, 16'hFFFF,
16'h12BB, 16'hFFFF,
16'h12BC, 16'hFFFF,
16'h12BD, 16'hFFFF,
16'h12BE, 16'hFFFF,
16'h12BF, 16'hFFFF,
16'h12C0, 16'hFFFF,
16'h12C1, 16'hFFFF,
16'h12C2, 16'hFFFF,
16'h12C3, 16'hFFFF,
16'h12C4, 16'hFFFF,
16'h12C5, 16'hFFFF,
16'h12C6, 16'hFFFF,
16'h12C7, 16'hFFFF,
16'h12C8, 16'hFFFF,
16'h12C9, 16'hFFFF,
16'h12CA, 16'hFFFF,
16'h12CB, 16'hFFFF,
16'h12CC, 16'hFFFF,
16'h12CD, 16'hFFFF,
16'h12CE, 16'hFFFF,
16'h12CF, 16'hFFFF,
16'h12D0, 16'hFFFF,
16'h12D1, 16'hFFFF,
16'h12D2, 16'hFFFF,
16'h12D3, 16'hFFFF,
16'h12D4, 16'hFFFF,
16'h12D5, 16'hFFFF,
16'h12D6, 16'hFFFF,
16'h12D7, 16'hFFFF,
16'h12D8, 16'hFFFF,
16'h12D9, 16'hFFFF,
16'h12DA, 16'hFFFF,
16'h12DB, 16'hFFFF,
16'h12DC, 16'hFFFF,
16'h12DD, 16'hFFFF,
16'h12DE, 16'hFFFF,
16'h12DF, 16'hFFFF,
16'h12E0, 16'hFFFF,
16'h12E1, 16'hFFFF,
16'h12E2, 16'hFFFF,
16'h12E3, 16'hFFFF,
16'h12E4, 16'hFFFF,
16'h12E5, 16'hFFFF,
16'h12E6, 16'hFFFF,
16'h12E7, 16'hFFFF,
16'h12E8, 16'hFFFF,
16'h12E9, 16'hFFFF,
16'h12EA, 16'hFFFF,
16'h12EB, 16'hFFFF,
16'h12EC, 16'hFFFF,
16'h12ED, 16'hFFFF,
16'h12EE, 16'hFFFF,
16'h12EF, 16'hFFFF,
16'h12F0, 16'hFFFF,
16'h12F1, 16'hFFFF,
16'h12F2, 16'hFFFF,
16'h12F3, 16'hFFFF,
16'h12F4, 16'hFFFF,
16'h12F5, 16'hFFFF,
16'h12F6, 16'hFFFF,
16'h12F7, 16'hFFFF,
16'h12F8, 16'hFFFF,
16'h12F9, 16'hFFFF,
16'h12FA, 16'hFFFF,
16'h12FB, 16'hFFFF,
16'h12FC, 16'hFFFF,
16'h12FD, 16'hFFFF,
16'h12FE, 16'hFFFF,
16'h12FF, 16'hFFFF,
16'h1300, 16'hFFFF,
16'h1301, 16'hFFFF,
16'h1302, 16'hFFFF,
16'h1303, 16'hFFFF,
16'h1304, 16'hFFFF,
16'h1305, 16'hFFFF,
16'h1306, 16'hFFFF,
16'h1307, 16'hFFFF,
16'h1308, 16'hFFFF,
16'h1309, 16'hFFFF,
16'h130A, 16'hFFFF,
16'h130B, 16'hFFFF,
16'h130C, 16'hFFFF,
16'h130D, 16'hFFFF,
16'h130E, 16'hFFFF,
16'h130F, 16'hFFFF,
16'h1310, 16'hFFFF,
16'h1311, 16'hFFFF,
16'h1312, 16'hFFFF,
16'h1313, 16'hFFFF,
16'h1314, 16'hFFFF,
16'h1315, 16'hFFFF,
16'h1316, 16'hFFFF,
16'h1317, 16'hFFFF,
16'h1318, 16'hFFFF,
16'h1319, 16'hFFFF,
16'h131A, 16'hFFFF,
16'h131B, 16'hFFFF,
16'h131C, 16'hFFFF,
16'h131D, 16'hFFFF,
16'h131E, 16'hFFFF,
16'h131F, 16'hFFFF,
16'h1320, 16'hFFFF,
16'h1321, 16'hFFFF,
16'h1322, 16'hFFFF,
16'h1323, 16'hFFFF,
16'h1324, 16'hFFFF,
16'h1325, 16'hFFFF,
16'h1326, 16'hFFFF,
16'h1327, 16'hFFFF,
16'h1328, 16'hFFFF,
16'h1329, 16'hFFFF,
16'h132A, 16'hFFFF,
16'h132B, 16'hFFFF,
16'h132C, 16'hFFFF,
16'h132D, 16'hFFFF,
16'h132E, 16'hFFFF,
16'h132F, 16'hFFFF,
16'h1330, 16'hFFFF,
16'h1331, 16'hFFFF,
16'h1332, 16'hFFFF,
16'h1333, 16'hFFFF,
16'h1334, 16'hFFFF,
16'h1335, 16'hFFFF,
16'h1336, 16'hFFFF,
16'h1337, 16'hFFFF,
16'h1338, 16'hFFFF,
16'h1339, 16'hFFFF,
16'h133A, 16'hFFFF,
16'h133B, 16'hFFFF,
16'h133C, 16'hFFFF,
16'h133D, 16'hFFFF,
16'h133E, 16'hFFFF,
16'h133F, 16'hFFFF,
16'h1340, 16'hFFFF,
16'h1341, 16'hFFFF,
16'h1342, 16'hFFFF,
16'h1343, 16'hFFFF,
16'h1344, 16'hFFFF,
16'h1345, 16'hFFFF,
16'h1346, 16'hFFFF,
16'h1347, 16'hFFFF,
16'h1348, 16'hFFFF,
16'h1349, 16'hFFFF,
16'h134A, 16'hFFFF,
16'h134B, 16'hFFFF,
16'h134C, 16'hFFFF,
16'h134D, 16'hFFFF,
16'h134E, 16'hFFFF,
16'h134F, 16'hFFFF,
16'h1350, 16'hFFFF,
16'h1351, 16'hFFFF,
16'h1352, 16'hFFFF,
16'h1353, 16'hFFFF,
16'h1354, 16'hFFFF,
16'h1355, 16'hFFFF,
16'h1356, 16'hFFFF,
16'h1357, 16'hFFFF,
16'h1358, 16'hFFFF,
16'h1359, 16'hFFFF,
16'h135A, 16'hFFFF,
16'h135B, 16'hFFFF,
16'h135C, 16'hFFFF,
16'h135D, 16'hFFFF,
16'h135E, 16'hFFFF,
16'h135F, 16'hFFFF,
16'h1360, 16'hFFFF,
16'h1361, 16'hFFFF,
16'h1362, 16'hFFFF,
16'h1363, 16'hFFFF,
16'h1364, 16'hFFFF,
16'h1365, 16'hFFFF,
16'h1366, 16'hFFFF,
16'h1367, 16'hFFFF,
16'h1368, 16'hFFFF,
16'h1369, 16'hFFFF,
16'h136A, 16'hFFFF,
16'h136B, 16'hFFFF,
16'h136C, 16'hFFFF,
16'h136D, 16'hFFFF,
16'h136E, 16'hFFFF,
16'h136F, 16'hFFFF,
16'h1370, 16'hFFFF,
16'h1371, 16'hFFFF,
16'h1372, 16'hFFFF,
16'h1373, 16'hFFFF,
16'h1374, 16'hFFFF,
16'h1375, 16'hFFFF,
16'h1376, 16'hFFFF,
16'h1377, 16'hFFFF,
16'h1378, 16'hFFFF,
16'h1379, 16'hFFFF,
16'h137A, 16'hFFFF,
16'h137B, 16'hFFFF,
16'h137C, 16'hFFFF,
16'h137D, 16'hFFFF,
16'h137E, 16'hFFFF,
16'h137F, 16'hFFFF,
16'h1380, 16'hFFFF,
16'h1381, 16'hFFFF,
16'h1382, 16'hFFFF,
16'h1383, 16'hFFFF,
16'h1384, 16'hFFFF,
16'h1385, 16'hFFFF,
16'h1386, 16'hFFFF,
16'h1387, 16'hFFFF,
16'h1388, 16'hFFFF,
16'h1389, 16'hFFFF,
16'h138A, 16'hFFFF,
16'h138B, 16'hFFFF,
16'h138C, 16'hFFFF,
16'h138D, 16'hFFFF,
16'h138E, 16'hFFFF,
16'h138F, 16'hFFFF,
16'h1390, 16'hFFFF,
16'h1391, 16'hFFFF,
16'h1392, 16'hFFFF,
16'h1393, 16'hFFFF,
16'h1394, 16'hFFFF,
16'h1395, 16'hFFFF,
16'h1396, 16'hFFFF,
16'h1397, 16'hFFFF,
16'h1398, 16'hFFFF,
16'h1399, 16'hFFFF,
16'h139A, 16'hFFFF,
16'h139B, 16'hFFFF,
16'h139C, 16'hFFFF,
16'h139D, 16'hFFFF,
16'h139E, 16'hFFFF,
16'h139F, 16'hFFFF,
16'h13A0, 16'hFFFF,
16'h13A1, 16'hFFFF,
16'h13A2, 16'hFFFF,
16'h13A3, 16'hFFFF,
16'h13A4, 16'hFFFF,
16'h13A5, 16'hFFFF,
16'h13A6, 16'hFFFF,
16'h13A7, 16'hFFFF,
16'h13A8, 16'hFFFF,
16'h13A9, 16'hFFFF,
16'h13AA, 16'hFFFF,
16'h13AB, 16'hFFFF,
16'h13AC, 16'hFFFF,
16'h13AD, 16'hFFFF,
16'h13AE, 16'hFFFF,
16'h13AF, 16'hFFFF,
16'h13B0, 16'hFFFF,
16'h13B1, 16'hFFFF,
16'h13B2, 16'hFFFF,
16'h13B3, 16'hFFFF,
16'h13B4, 16'hFFFF,
16'h13B5, 16'hFFFF,
16'h13B6, 16'hFFFF,
16'h13B7, 16'hFFFF,
16'h13B8, 16'hFFFF,
16'h13B9, 16'hFFFF,
16'h13BA, 16'hFFFF,
16'h13BB, 16'hFFFF,
16'h13BC, 16'hFFFF,
16'h13BD, 16'hFFFF,
16'h13BE, 16'hFFFF,
16'h13BF, 16'hFFFF,
16'h13C0, 16'hFFFF,
16'h13C1, 16'hFFFF,
16'h13C2, 16'hFFFF,
16'h13C3, 16'hFFFF,
16'h13C4, 16'hFFFF,
16'h13C5, 16'hFFFF,
16'h13C6, 16'hFFFF,
16'h13C7, 16'hFFFF,
16'h13C8, 16'hFFFF,
16'h13C9, 16'hFFFF,
16'h13CA, 16'hFFFF,
16'h13CB, 16'hFFFF,
16'h13CC, 16'hFFFF,
16'h13CD, 16'hFFFF,
16'h13CE, 16'hFFFF,
16'h13CF, 16'hFFFF,
16'h13D0, 16'hFFFF,
16'h13D1, 16'hFFFF,
16'h13D2, 16'hFFFF,
16'h13D3, 16'hFFFF,
16'h13D4, 16'hFFFF,
16'h13D5, 16'hFFFF,
16'h13D6, 16'hFFFF,
16'h13D7, 16'hFFFF,
16'h13D8, 16'hFFFF,
16'h13D9, 16'hFFFF,
16'h13DA, 16'hFFFF,
16'h13DB, 16'hFFFF,
16'h13DC, 16'hFFFF,
16'h13DD, 16'hFFFF,
16'h13DE, 16'hFFFF,
16'h13DF, 16'hFFFF,
16'h13E0, 16'hFFFF,
16'h13E1, 16'hFFFF,
16'h13E2, 16'hFFFF,
16'h13E3, 16'hFFFF,
16'h13E4, 16'hFFFF,
16'h13E5, 16'hFFFF,
16'h13E6, 16'hFFFF,
16'h13E7, 16'hFFFF,
16'h13E8, 16'hFFFF,
16'h13E9, 16'hFFFF,
16'h13EA, 16'hFFFF,
16'h13EB, 16'hFFFF,
16'h13EC, 16'hFFFF,
16'h13ED, 16'hFFFF,
16'h13EE, 16'hFFFF,
16'h13EF, 16'hFFFF,
16'h13F0, 16'hFFFF,
16'h13F1, 16'hFFFF,
16'h13F2, 16'hFFFF,
16'h13F3, 16'hFFFF,
16'h13F4, 16'hFFFF,
16'h13F5, 16'hFFFF,
16'h13F6, 16'hFFFF,
16'h13F7, 16'hFFFF,
16'h13F8, 16'hFFFF,
16'h13F9, 16'hFFFF,
16'h13FA, 16'hFFFF,
16'h13FB, 16'hFFFF,
16'h13FC, 16'hFFFF,
16'h13FD, 16'hFFFF,
16'h13FE, 16'hFFFF,
16'h13FF, 16'hFFFF,
16'h1400, 16'hFFFF,
16'h1401, 16'hFFFF,
16'h1402, 16'hFFFF,
16'h1403, 16'hFFFF,
16'h1404, 16'hFFFF,
16'h1405, 16'hFFFF,
16'h1406, 16'hFFFF,
16'h1407, 16'hFFFF,
16'h1408, 16'hFFFF,
16'h1409, 16'hFFFF,
16'h140A, 16'hFFFF,
16'h140B, 16'hFFFF,
16'h140C, 16'hFFFF,
16'h140D, 16'hFFFF,
16'h140E, 16'hFFFF,
16'h140F, 16'hFFFF,
16'h1410, 16'hFFFF,
16'h1411, 16'hFFFF,
16'h1412, 16'hFFFF,
16'h1413, 16'hFFFF,
16'h1414, 16'hFFFF,
16'h1415, 16'hFFFF,
16'h1416, 16'hFFFF,
16'h1417, 16'hFFFF,
16'h1418, 16'hFFFF,
16'h1419, 16'hFFFF,
16'h141A, 16'hFFFF,
16'h141B, 16'hFFFF,
16'h141C, 16'hFFFF,
16'h141D, 16'hFFFF,
16'h141E, 16'hFFFF,
16'h141F, 16'hFFFF,
16'h1420, 16'hFFFF,
16'h1421, 16'hFFFF,
16'h1422, 16'hFFFF,
16'h1423, 16'hFFFF,
16'h1424, 16'hFFFF,
16'h1425, 16'hFFFF,
16'h1426, 16'hFFFF,
16'h1427, 16'hFFFF,
16'h1428, 16'hFFFF,
16'h1429, 16'hFFFF,
16'h142A, 16'hFFFF,
16'h142B, 16'hFFFF,
16'h142C, 16'hFFFF,
16'h142D, 16'hFFFF,
16'h142E, 16'hFFFF,
16'h142F, 16'hFFFF,
16'h1430, 16'hFFFF,
16'h1431, 16'hFFFF,
16'h1432, 16'hFFFF,
16'h1433, 16'hFFFF,
16'h1434, 16'hFFFF,
16'h1435, 16'hFFFF,
16'h1436, 16'hFFFF,
16'h1437, 16'hFFFF,
16'h1438, 16'hFFFF,
16'h1439, 16'hFFFF,
16'h143A, 16'hFFFF,
16'h143B, 16'hFFFF,
16'h143C, 16'hFFFF,
16'h143D, 16'hFFFF,
16'h143E, 16'hFFFF,
16'h143F, 16'hFFFF,
16'h1440, 16'hFFFF,
16'h1441, 16'hFFFF,
16'h1442, 16'hFFFF,
16'h1443, 16'hFFFF,
16'h1444, 16'hFFFF,
16'h1445, 16'hFFFF,
16'h1446, 16'hFFFF,
16'h1447, 16'hFFFF,
16'h1448, 16'hFFFF,
16'h1449, 16'hFFFF,
16'h144A, 16'hFFFF,
16'h144B, 16'hFFFF,
16'h144C, 16'hFFFF,
16'h144D, 16'hFFFF,
16'h144E, 16'hFFFF,
16'h144F, 16'hFFFF,
16'h1450, 16'hFFFF,
16'h1451, 16'hFFFF,
16'h1452, 16'hFFFF,
16'h1453, 16'hFFFF,
16'h1454, 16'hFFFF,
16'h1455, 16'hFFFF,
16'h1456, 16'hFFFF,
16'h1457, 16'hFFFF,
16'h1458, 16'hFFFF,
16'h1459, 16'hFFFF,
16'h145A, 16'hFFFF,
16'h145B, 16'hFFFF,
16'h145C, 16'hFFFF,
16'h145D, 16'hFFFF,
16'h145E, 16'hFFFF,
16'h145F, 16'hFFFF,
16'h1460, 16'hFFFF,
16'h1461, 16'hFFFF,
16'h1462, 16'hFFFF,
16'h1463, 16'hFFFF,
16'h1464, 16'hFFFF,
16'h1465, 16'hFFFF,
16'h1466, 16'hFFFF,
16'h1467, 16'hFFFF,
16'h1468, 16'hFFFF,
16'h1469, 16'hFFFF,
16'h146A, 16'hFFFF,
16'h146B, 16'hFFFF,
16'h146C, 16'hFFFF,
16'h146D, 16'hFFFF,
16'h146E, 16'hFFFF,
16'h146F, 16'hFFFF,
16'h1470, 16'hFFFF,
16'h1471, 16'hFFFF,
16'h1472, 16'hFFFF,
16'h1473, 16'hFFFF,
16'h1474, 16'hFFFF,
16'h1475, 16'hFFFF,
16'h1476, 16'hFFFF,
16'h1477, 16'hFFFF,
16'h1478, 16'hFFFF,
16'h1479, 16'hFFFF,
16'h147A, 16'hFFFF,
16'h147B, 16'hFFFF,
16'h147C, 16'hFFFF,
16'h147D, 16'hFFFF,
16'h147E, 16'hFFFF,
16'h147F, 16'hFFFF,
16'h1480, 16'hFFFF,
16'h1481, 16'hFFFF,
16'h1482, 16'hFFFF,
16'h1483, 16'hFFFF,
16'h1484, 16'hFFFF,
16'h1485, 16'hFFFF,
16'h1486, 16'hFFFF,
16'h1487, 16'hFFFF,
16'h1488, 16'hFFFF,
16'h1489, 16'hFFFF,
16'h148A, 16'hFFFF,
16'h148B, 16'hFFFF,
16'h148C, 16'hFFFF,
16'h148D, 16'hFFFF,
16'h148E, 16'hFFFF,
16'h148F, 16'hFFFF,
16'h1490, 16'hFFFF,
16'h1491, 16'hFFFF,
16'h1492, 16'hFFFF,
16'h1493, 16'hFFFF,
16'h1494, 16'hFFFF,
16'h1495, 16'hFFFF,
16'h1496, 16'hFFFF,
16'h1497, 16'hFFFF,
16'h1498, 16'hFFFF,
16'h1499, 16'hFFFF,
16'h149A, 16'hFFFF,
16'h149B, 16'hFFFF,
16'h149C, 16'hFFFF,
16'h149D, 16'hFFFF,
16'h149E, 16'hFFFF,
16'h149F, 16'hFFFF,
16'h14A0, 16'hFFFF,
16'h14A1, 16'hFFFF,
16'h14A2, 16'hFFFF,
16'h14A3, 16'hFFFF,
16'h14A4, 16'hFFFF,
16'h14A5, 16'hFFFF,
16'h14A6, 16'hFFFF,
16'h14A7, 16'hFFFF,
16'h14A8, 16'hFFFF,
16'h14A9, 16'hFFFF,
16'h14AA, 16'hFFFF,
16'h14AB, 16'hFFFF,
16'h14AC, 16'hFFFF,
16'h14AD, 16'hFFFF,
16'h14AE, 16'hFFFF,
16'h14AF, 16'hFFFF,
16'h14B0, 16'hFFFF,
16'h14B1, 16'hFFFF,
16'h14B2, 16'hFFFF,
16'h14B3, 16'hFFFF,
16'h14B4, 16'hFFFF,
16'h14B5, 16'hFFFF,
16'h14B6, 16'hFFFF,
16'h14B7, 16'hFFFF,
16'h14B8, 16'hFFFF,
16'h14B9, 16'hFFFF,
16'h14BA, 16'hFFFF,
16'h14BB, 16'hFFFF,
16'h14BC, 16'hFFFF,
16'h14BD, 16'hFFFF,
16'h14BE, 16'hFFFF,
16'h14BF, 16'hFFFF,
16'h14C0, 16'hFFFF,
16'h14C1, 16'hFFFF,
16'h14C2, 16'hFFFF,
16'h14C3, 16'hFFFF,
16'h14C4, 16'hFFFF,
16'h14C5, 16'hFFFF,
16'h14C6, 16'hFFFF,
16'h14C7, 16'hFFFF,
16'h14C8, 16'hFFFF,
16'h14C9, 16'hFFFF,
16'h14CA, 16'hFFFF,
16'h14CB, 16'hFFFF,
16'h14CC, 16'hFFFF,
16'h14CD, 16'hFFFF,
16'h14CE, 16'hFFFF,
16'h14CF, 16'hFFFF,
16'h14D0, 16'hFFFF,
16'h14D1, 16'hFFFF,
16'h14D2, 16'hFFFF,
16'h14D3, 16'hFFFF,
16'h14D4, 16'hFFFF,
16'h14D5, 16'hFFFF,
16'h14D6, 16'hFFFF,
16'h14D7, 16'hFFFF,
16'h14D8, 16'hFFFF,
16'h14D9, 16'hFFFF,
16'h14DA, 16'hFFFF,
16'h14DB, 16'hFFFF,
16'h14DC, 16'hFFFF,
16'h14DD, 16'hFFFF,
16'h14DE, 16'hFFFF,
16'h14DF, 16'hFFFF,
16'h14E0, 16'hFFFF,
16'h14E1, 16'hFFFF,
16'h14E2, 16'hFFFF,
16'h14E3, 16'hFFFF,
16'h14E4, 16'hFFFF,
16'h14E5, 16'hFFFF,
16'h14E6, 16'hFFFF,
16'h14E7, 16'hFFFF,
16'h14E8, 16'hFFFF,
16'h14E9, 16'hFFFF,
16'h14EA, 16'hFFFF,
16'h14EB, 16'hFFFF,
16'h14EC, 16'hFFFF,
16'h14ED, 16'hFFFF,
16'h14EE, 16'hFFFF,
16'h14EF, 16'hFFFF,
16'h14F0, 16'hFFFF,
16'h14F1, 16'hFFFF,
16'h14F2, 16'hFFFF,
16'h14F3, 16'hFFFF,
16'h14F4, 16'hFFFF,
16'h14F5, 16'hFFFF,
16'h14F6, 16'hFFFF,
16'h14F7, 16'hFFFF,
16'h14F8, 16'hFFFF,
16'h14F9, 16'hFFFF,
16'h14FA, 16'hFFFF,
16'h14FB, 16'hFFFF,
16'h14FC, 16'hFFFF,
16'h14FD, 16'hFFFF,
16'h14FE, 16'hFFFF,
16'h14FF, 16'hFFFF,
16'h1500, 16'hFFFF,
16'h1501, 16'hFFFF,
16'h1502, 16'hFFFF,
16'h1503, 16'hFFFF,
16'h1504, 16'hFFFF,
16'h1505, 16'hFFFF,
16'h1506, 16'hFFFF,
16'h1507, 16'hFFFF,
16'h1508, 16'hFFFF,
16'h1509, 16'hFFFF,
16'h150A, 16'hFFFF,
16'h150B, 16'hFFFF,
16'h150C, 16'hFFFF,
16'h150D, 16'hFFFF,
16'h150E, 16'hFFFF,
16'h150F, 16'hFFFF,
16'h1510, 16'hFFFF,
16'h1511, 16'hFFFF,
16'h1512, 16'hFFFF,
16'h1513, 16'hFFFF,
16'h1514, 16'hFFFF,
16'h1515, 16'hFFFF,
16'h1516, 16'hFFFF,
16'h1517, 16'hFFFF,
16'h1518, 16'hFFFF,
16'h1519, 16'hFFFF,
16'h151A, 16'hFFFF,
16'h151B, 16'hFFFF,
16'h151C, 16'hFFFF,
16'h151D, 16'hFFFF,
16'h151E, 16'hFFFF,
16'h151F, 16'hFFFF,
16'h1520, 16'hFFFF,
16'h1521, 16'hFFFF,
16'h1522, 16'hFFFF,
16'h1523, 16'hFFFF,
16'h1524, 16'hFFFF,
16'h1525, 16'hFFFF,
16'h1526, 16'hFFFF,
16'h1527, 16'hFFFF,
16'h1528, 16'hFFFF,
16'h1529, 16'hFFFF,
16'h152A, 16'hFFFF,
16'h152B, 16'hFFFF,
16'h152C, 16'hFFFF,
16'h152D, 16'hFFFF,
16'h152E, 16'hFFFF,
16'h152F, 16'hFFFF,
16'h1530, 16'hFFFF,
16'h1531, 16'hFFFF,
16'h1532, 16'hFFFF,
16'h1533, 16'hFFFF,
16'h1534, 16'hFFFF,
16'h1535, 16'hFFFF,
16'h1536, 16'hFFFF,
16'h1537, 16'hFFFF,
16'h1538, 16'hFFFF,
16'h1539, 16'hFFFF,
16'h153A, 16'hFFFF,
16'h153B, 16'hFFFF,
16'h153C, 16'hFFFF,
16'h153D, 16'hFFFF,
16'h153E, 16'hFFFF,
16'h153F, 16'hFFFF,
16'h1540, 16'hFFFF,
16'h1541, 16'hFFFF,
16'h1542, 16'hFFFF,
16'h1543, 16'hFFFF,
16'h1544, 16'hFFFF,
16'h1545, 16'hFFFF,
16'h1546, 16'hFFFF,
16'h1547, 16'hFFFF,
16'h1548, 16'hFFFF,
16'h1549, 16'hFFFF,
16'h154A, 16'hFFFF,
16'h154B, 16'hFFFF,
16'h154C, 16'hFFFF,
16'h154D, 16'hFFFF,
16'h154E, 16'hFFFF,
16'h154F, 16'hFFFF,
16'h1550, 16'hFFFF,
16'h1551, 16'hFFFF,
16'h1552, 16'hFFFF,
16'h1553, 16'hFFFF,
16'h1554, 16'hFFFF,
16'h1555, 16'hFFFF,
16'h1556, 16'hFFFF,
16'h1557, 16'hFFFF,
16'h1558, 16'hFFFF,
16'h1559, 16'hFFFF,
16'h155A, 16'hFFFF,
16'h155B, 16'hFFFF,
16'h155C, 16'hFFFF,
16'h155D, 16'hFFFF,
16'h155E, 16'hFFFF,
16'h155F, 16'hFFFF,
16'h1560, 16'hFFFF,
16'h1561, 16'hFFFF,
16'h1562, 16'hFFFF,
16'h1563, 16'hFFFF,
16'h1564, 16'hFFFF,
16'h1565, 16'hFFFF,
16'h1566, 16'hFFFF,
16'h1567, 16'hFFFF,
16'h1568, 16'hFFFF,
16'h1569, 16'hFFFF,
16'h156A, 16'hFFFF,
16'h156B, 16'hFFFF,
16'h156C, 16'hFFFF,
16'h156D, 16'hFFFF,
16'h156E, 16'hFFFF,
16'h156F, 16'hFFFF,
16'h1570, 16'hFFFF,
16'h1571, 16'hFFFF,
16'h1572, 16'hFFFF,
16'h1573, 16'hFFFF,
16'h1574, 16'hFFFF,
16'h1575, 16'hFFFF,
16'h1576, 16'hFFFF,
16'h1577, 16'hFFFF,
16'h1578, 16'hFFFF,
16'h1579, 16'hFFFF,
16'h157A, 16'hFFFF,
16'h157B, 16'hFFFF,
16'h157C, 16'hFFFF,
16'h157D, 16'hFFFF,
16'h157E, 16'hFFFF,
16'h157F, 16'hFFFF,
16'h1580, 16'hFFFF,
16'h1581, 16'hFFFF,
16'h1582, 16'hFFFF,
16'h1583, 16'hFFFF,
16'h1584, 16'hFFFF,
16'h1585, 16'hFFFF,
16'h1586, 16'hFFFF,
16'h1587, 16'hFFFF,
16'h1588, 16'hFFFF,
16'h1589, 16'hFFFF,
16'h158A, 16'hFFFF,
16'h158B, 16'hFFFF,
16'h158C, 16'hFFFF,
16'h158D, 16'hFFFF,
16'h158E, 16'hFFFF,
16'h158F, 16'hFFFF,
16'h1590, 16'hFFFF,
16'h1591, 16'hFFFF,
16'h1592, 16'hFFFF,
16'h1593, 16'hFFFF,
16'h1594, 16'hFFFF,
16'h1595, 16'hFFFF,
16'h1596, 16'hFFFF,
16'h1597, 16'hFFFF,
16'h1598, 16'hFFFF,
16'h1599, 16'hFFFF,
16'h159A, 16'hFFFF,
16'h159B, 16'hFFFF,
16'h159C, 16'hFFFF,
16'h159D, 16'hFFFF,
16'h159E, 16'hFFFF,
16'h159F, 16'hFFFF,
16'h15A0, 16'hFFFF,
16'h15A1, 16'hFFFF,
16'h15A2, 16'hFFFF,
16'h15A3, 16'hFFFF,
16'h15A4, 16'hFFFF,
16'h15A5, 16'hFFFF,
16'h15A6, 16'hFFFF,
16'h15A7, 16'hFFFF,
16'h15A8, 16'hFFFF,
16'h15A9, 16'hFFFF,
16'h15AA, 16'hFFFF,
16'h15AB, 16'hFFFF,
16'h15AC, 16'hFFFF,
16'h15AD, 16'hFFFF,
16'h15AE, 16'hFFFF,
16'h15AF, 16'hFFFF,
16'h15B0, 16'hFFFF,
16'h15B1, 16'hFFFF,
16'h15B2, 16'hFFFF,
16'h15B3, 16'hFFFF,
16'h15B4, 16'hFFFF,
16'h15B5, 16'hFFFF,
16'h15B6, 16'hFFFF,
16'h15B7, 16'hFFFF,
16'h15B8, 16'hFFFF,
16'h15B9, 16'hFFFF,
16'h15BA, 16'hFFFF,
16'h15BB, 16'hFFFF,
16'h15BC, 16'hFFFF,
16'h15BD, 16'hFFFF,
16'h15BE, 16'hFFFF,
16'h15BF, 16'hFFFF,
16'h15C0, 16'hFFFF,
16'h15C1, 16'hFFFF,
16'h15C2, 16'hFFFF,
16'h15C3, 16'hFFFF,
16'h15C4, 16'hFFFF,
16'h15C5, 16'hFFFF,
16'h15C6, 16'hFFFF,
16'h15C7, 16'hFFFF,
16'h15C8, 16'hFFFF,
16'h15C9, 16'hFFFF,
16'h15CA, 16'hFFFF,
16'h15CB, 16'hFFFF,
16'h15CC, 16'hFFFF,
16'h15CD, 16'hFFFF,
16'h15CE, 16'hFFFF,
16'h15CF, 16'hFFFF,
16'h15D0, 16'hFFFF,
16'h15D1, 16'hFFFF,
16'h15D2, 16'hFFFF,
16'h15D3, 16'hFFFF,
16'h15D4, 16'hFFFF,
16'h15D5, 16'hFFFF,
16'h15D6, 16'hFFFF,
16'h15D7, 16'hFFFF,
16'h15D8, 16'hFFFF,
16'h15D9, 16'hFFFF,
16'h15DA, 16'hFFFF,
16'h15DB, 16'hFFFF,
16'h15DC, 16'hFFFF,
16'h15DD, 16'hFFFF,
16'h15DE, 16'hFFFF,
16'h15DF, 16'hFFFF,
16'h15E0, 16'hFFFF,
16'h15E1, 16'hFFFF,
16'h15E2, 16'hFFFF,
16'h15E3, 16'hFFFF,
16'h15E4, 16'hFFFF,
16'h15E5, 16'hFFFF,
16'h15E6, 16'hFFFF,
16'h15E7, 16'hFFFF,
16'h15E8, 16'hFFFF,
16'h15E9, 16'hFFFF,
16'h15EA, 16'hFFFF,
16'h15EB, 16'hFFFF,
16'h15EC, 16'hFFFF,
16'h15ED, 16'hFFFF,
16'h15EE, 16'hFFFF,
16'h15EF, 16'hFFFF,
16'h15F0, 16'hFFFF,
16'h15F1, 16'hFFFF,
16'h15F2, 16'hFFFF,
16'h15F3, 16'hFFFF,
16'h15F4, 16'hFFFF,
16'h15F5, 16'hFFFF,
16'h15F6, 16'hFFFF,
16'h15F7, 16'hFFFF,
16'h15F8, 16'hFFFF,
16'h15F9, 16'hFFFF,
16'h15FA, 16'hFFFF,
16'h15FB, 16'hFFFF,
16'h15FC, 16'hFFFF,
16'h15FD, 16'hFFFF,
16'h15FE, 16'hFFFF,
16'h15FF, 16'hFFFF,
16'h1600, 16'hFFFF,
16'h1601, 16'hFFFF,
16'h1602, 16'hFFFF,
16'h1603, 16'hFFFF,
16'h1604, 16'hFFFF,
16'h1605, 16'hFFFF,
16'h1606, 16'hFFFF,
16'h1607, 16'hFFFF,
16'h1608, 16'hFFFF,
16'h1609, 16'hFFFF,
16'h160A, 16'hFFFF,
16'h160B, 16'hFFFF,
16'h160C, 16'hFFFF,
16'h160D, 16'hFFFF,
16'h160E, 16'hFFFF,
16'h160F, 16'hFFFF,
16'h1610, 16'hFFFF,
16'h1611, 16'hFFFF,
16'h1612, 16'hFFFF,
16'h1613, 16'hFFFF,
16'h1614, 16'hFFFF,
16'h1615, 16'hFFFF,
16'h1616, 16'hFFFF,
16'h1617, 16'hFFFF,
16'h1618, 16'hFFFF,
16'h1619, 16'hFFFF,
16'h161A, 16'hFFFF,
16'h161B, 16'hFFFF,
16'h161C, 16'hFFFF,
16'h161D, 16'hFFFF,
16'h161E, 16'hFFFF,
16'h161F, 16'hFFFF,
16'h1620, 16'hFFFF,
16'h1621, 16'hFFFF,
16'h1622, 16'hFFFF,
16'h1623, 16'hFFFF,
16'h1624, 16'hFFFF,
16'h1625, 16'hFFFF,
16'h1626, 16'hFFFF,
16'h1627, 16'hFFFF,
16'h1628, 16'hFFFF,
16'h1629, 16'hFFFF,
16'h162A, 16'hFFFF,
16'h162B, 16'hFFFF,
16'h162C, 16'hFFFF,
16'h162D, 16'hFFFF,
16'h162E, 16'hFFFF,
16'h162F, 16'hFFFF,
16'h1630, 16'hFFFF,
16'h1631, 16'hFFFF,
16'h1632, 16'hFFFF,
16'h1633, 16'hFFFF,
16'h1634, 16'hFFFF,
16'h1635, 16'hFFFF,
16'h1636, 16'hFFFF,
16'h1637, 16'hFFFF,
16'h1638, 16'hFFFF,
16'h1639, 16'hFFFF,
16'h163A, 16'hFFFF,
16'h163B, 16'hFFFF,
16'h163C, 16'hFFFF,
16'h163D, 16'hFFFF,
16'h163E, 16'hFFFF,
16'h163F, 16'hFFFF,
16'h1640, 16'hFFFF,
16'h1641, 16'hFFFF,
16'h1642, 16'hFFFF,
16'h1643, 16'hFFFF,
16'h1644, 16'hFFFF,
16'h1645, 16'hFFFF,
16'h1646, 16'hFFFF,
16'h1647, 16'hFFFF,
16'h1648, 16'hFFFF,
16'h1649, 16'hFFFF,
16'h164A, 16'hFFFF,
16'h164B, 16'hFFFF,
16'h164C, 16'hFFFF,
16'h164D, 16'hFFFF,
16'h164E, 16'hFFFF,
16'h164F, 16'hFFFF,
16'h1650, 16'hFFFF,
16'h1651, 16'hFFFF,
16'h1652, 16'hFFFF,
16'h1653, 16'hFFFF,
16'h1654, 16'hFFFF,
16'h1655, 16'hFFFF,
16'h1656, 16'hFFFF,
16'h1657, 16'hFFFF,
16'h1658, 16'hFFFF,
16'h1659, 16'hFFFF,
16'h165A, 16'hFFFF,
16'h165B, 16'hFFFF,
16'h165C, 16'hFFFF,
16'h165D, 16'hFFFF,
16'h165E, 16'hFFFF,
16'h165F, 16'hFFFF,
16'h1660, 16'hFFFF,
16'h1661, 16'hFFFF,
16'h1662, 16'hFFFF,
16'h1663, 16'hFFFF,
16'h1664, 16'hFFFF,
16'h1665, 16'hFFFF,
16'h1666, 16'hFFFF,
16'h1667, 16'hFFFF,
16'h1668, 16'hFFFF,
16'h1669, 16'hFFFF,
16'h166A, 16'hFFFF,
16'h166B, 16'hFFFF,
16'h166C, 16'hFFFF,
16'h166D, 16'hFFFF,
16'h166E, 16'hFFFF,
16'h166F, 16'hFFFF,
16'h1670, 16'hFFFF,
16'h1671, 16'hFFFF,
16'h1672, 16'hFFFF,
16'h1673, 16'hFFFF,
16'h1674, 16'hFFFF,
16'h1675, 16'hFFFF,
16'h1676, 16'hFFFF,
16'h1677, 16'hFFFF,
16'h1678, 16'hFFFF,
16'h1679, 16'hFFFF,
16'h167A, 16'hFFFF,
16'h167B, 16'hFFFF,
16'h167C, 16'hFFFF,
16'h167D, 16'hFFFF,
16'h167E, 16'hFFFF,
16'h167F, 16'hFFFF,
16'h1680, 16'hFFFF,
16'h1681, 16'hFFFF,
16'h1682, 16'hFFFF,
16'h1683, 16'hFFFF,
16'h1684, 16'hFFFF,
16'h1685, 16'hFFFF,
16'h1686, 16'hFFFF,
16'h1687, 16'hFFFF,
16'h1688, 16'hFFFF,
16'h1689, 16'hFFFF,
16'h168A, 16'hFFFF,
16'h168B, 16'hFFFF,
16'h168C, 16'hFFFF,
16'h168D, 16'hFFFF,
16'h168E, 16'hFFFF,
16'h168F, 16'hFFFF,
16'h1690, 16'hFFFF,
16'h1691, 16'hFFFF,
16'h1692, 16'hFFFF,
16'h1693, 16'hFFFF,
16'h1694, 16'hFFFF,
16'h1695, 16'hFFFF,
16'h1696, 16'hFFFF,
16'h1697, 16'hFFFF,
16'h1698, 16'hFFFF,
16'h1699, 16'hFFFF,
16'h169A, 16'hFFFF,
16'h169B, 16'hFFFF,
16'h169C, 16'hFFFF,
16'h169D, 16'hFFFF,
16'h169E, 16'hFFFF,
16'h169F, 16'hFFFF,
16'h16A0, 16'hFFFF,
16'h16A1, 16'hFFFF,
16'h16A2, 16'hFFFF,
16'h16A3, 16'hFFFF,
16'h16A4, 16'hFFFF,
16'h16A5, 16'hFFFF,
16'h16A6, 16'hFFFF,
16'h16A7, 16'hFFFF,
16'h16A8, 16'hFFFF,
16'h16A9, 16'hFFFF,
16'h16AA, 16'hFFFF,
16'h16AB, 16'hFFFF,
16'h16AC, 16'hFFFF,
16'h16AD, 16'hFFFF,
16'h16AE, 16'hFFFF,
16'h16AF, 16'hFFFF,
16'h16B0, 16'hFFFF,
16'h16B1, 16'hFFFF,
16'h16B2, 16'hFFFF,
16'h16B3, 16'hFFFF,
16'h16B4, 16'hFFFF,
16'h16B5, 16'hFFFF,
16'h16B6, 16'hFFFF,
16'h16B7, 16'hFFFF,
16'h16B8, 16'hFFFF,
16'h16B9, 16'hFFFF,
16'h16BA, 16'hFFFF,
16'h16BB, 16'hFFFF,
16'h16BC, 16'hFFFF,
16'h16BD, 16'hFFFF,
16'h16BE, 16'hFFFF,
16'h16BF, 16'hFFFF,
16'h16C0, 16'hFFFF,
16'h16C1, 16'hFFFF,
16'h16C2, 16'hFFFF,
16'h16C3, 16'hFFFF,
16'h16C4, 16'hFFFF,
16'h16C5, 16'hFFFF,
16'h16C6, 16'hFFFF,
16'h16C7, 16'hFFFF,
16'h16C8, 16'hFFFF,
16'h16C9, 16'hFFFF,
16'h16CA, 16'hFFFF,
16'h16CB, 16'hFFFF,
16'h16CC, 16'hFFFF,
16'h16CD, 16'hFFFF,
16'h16CE, 16'hFFFF,
16'h16CF, 16'hFFFF,
16'h16D0, 16'hFFFF,
16'h16D1, 16'hFFFF,
16'h16D2, 16'hFFFF,
16'h16D3, 16'hFFFF,
16'h16D4, 16'hFFFF,
16'h16D5, 16'hFFFF,
16'h16D6, 16'hFFFF,
16'h16D7, 16'hFFFF,
16'h16D8, 16'hFFFF,
16'h16D9, 16'hFFFF,
16'h16DA, 16'hFFFF,
16'h16DB, 16'hFFFF,
16'h16DC, 16'hFFFF,
16'h16DD, 16'hFFFF,
16'h16DE, 16'hFFFF,
16'h16DF, 16'hFFFF,
16'h16E0, 16'hFFFF,
16'h16E1, 16'hFFFF,
16'h16E2, 16'hFFFF,
16'h16E3, 16'hFFFF,
16'h16E4, 16'hFFFF,
16'h16E5, 16'hFFFF,
16'h16E6, 16'hFFFF,
16'h16E7, 16'hFFFF,
16'h16E8, 16'hFFFF,
16'h16E9, 16'hFFFF,
16'h16EA, 16'hFFFF,
16'h16EB, 16'hFFFF,
16'h16EC, 16'hFFFF,
16'h16ED, 16'hFFFF,
16'h16EE, 16'hFFFF,
16'h16EF, 16'hFFFF,
16'h16F0, 16'hFFFF,
16'h16F1, 16'hFFFF,
16'h16F2, 16'hFFFF,
16'h16F3, 16'hFFFF,
16'h16F4, 16'hFFFF,
16'h16F5, 16'hFFFF,
16'h16F6, 16'hFFFF,
16'h16F7, 16'hFFFF,
16'h16F8, 16'hFFFF,
16'h16F9, 16'hFFFF,
16'h16FA, 16'hFFFF,
16'h16FB, 16'hFFFF,
16'h16FC, 16'hFFFF,
16'h16FD, 16'hFFFF,
16'h16FE, 16'hFFFF,
16'h16FF, 16'hFFFF,
16'h1700, 16'hFFFF,
16'h1701, 16'hFFFF,
16'h1702, 16'hFFFF,
16'h1703, 16'hFFFF,
16'h1704, 16'hFFFF,
16'h1705, 16'hFFFF,
16'h1706, 16'hFFFF,
16'h1707, 16'hFFFF,
16'h1708, 16'hFFFF,
16'h1709, 16'hFFFF,
16'h170A, 16'hFFFF,
16'h170B, 16'hFFFF,
16'h170C, 16'hFFFF,
16'h170D, 16'hFFFF,
16'h170E, 16'hFFFF,
16'h170F, 16'hFFFF,
16'h1710, 16'hFFFF,
16'h1711, 16'hFFFF,
16'h1712, 16'hFFFF,
16'h1713, 16'hFFFF,
16'h1714, 16'hFFFF,
16'h1715, 16'hFFFF,
16'h1716, 16'hFFFF,
16'h1717, 16'hFFFF,
16'h1718, 16'hFFFF,
16'h1719, 16'hFFFF,
16'h171A, 16'hFFFF,
16'h171B, 16'hFFFF,
16'h171C, 16'hFFFF,
16'h171D, 16'hFFFF,
16'h171E, 16'hFFFF,
16'h171F, 16'hFFFF,
16'h1720, 16'hFFFF,
16'h1721, 16'hFFFF,
16'h1722, 16'hFFFF,
16'h1723, 16'hFFFF,
16'h1724, 16'hFFFF,
16'h1725, 16'hFFFF,
16'h1726, 16'hFFFF,
16'h1727, 16'hFFFF,
16'h1728, 16'hFFFF,
16'h1729, 16'hFFFF,
16'h172A, 16'hFFFF,
16'h172B, 16'hFFFF,
16'h172C, 16'hFFFF,
16'h172D, 16'hFFFF,
16'h172E, 16'hFFFF,
16'h172F, 16'hFFFF,
16'h1730, 16'hFFFF,
16'h1731, 16'hFFFF,
16'h1732, 16'hFFFF,
16'h1733, 16'hFFFF,
16'h1734, 16'hFFFF,
16'h1735, 16'hFFFF,
16'h1736, 16'hFFFF,
16'h1737, 16'hFFFF,
16'h1738, 16'hFFFF,
16'h1739, 16'hFFFF,
16'h173A, 16'hFFFF,
16'h173B, 16'hFFFF,
16'h173C, 16'hFFFF,
16'h173D, 16'hFFFF,
16'h173E, 16'hFFFF,
16'h173F, 16'hFFFF,
16'h1740, 16'hFFFF,
16'h1741, 16'hFFFF,
16'h1742, 16'hFFFF,
16'h1743, 16'hFFFF,
16'h1744, 16'hFFFF,
16'h1745, 16'hFFFF,
16'h1746, 16'hFFFF,
16'h1747, 16'hFFFF,
16'h1748, 16'hFFFF,
16'h1749, 16'hFFFF,
16'h174A, 16'hFFFF,
16'h174B, 16'hFFFF,
16'h174C, 16'hFFFF,
16'h174D, 16'hFFFF,
16'h174E, 16'hFFFF,
16'h174F, 16'hFFFF,
16'h1750, 16'hFFFF,
16'h1751, 16'hFFFF,
16'h1752, 16'hFFFF,
16'h1753, 16'hFFFF,
16'h1754, 16'hFFFF,
16'h1755, 16'hFFFF,
16'h1756, 16'hFFFF,
16'h1757, 16'hFFFF,
16'h1758, 16'hFFFF,
16'h1759, 16'hFFFF,
16'h175A, 16'hFFFF,
16'h175B, 16'hFFFF,
16'h175C, 16'hFFFF,
16'h175D, 16'hFFFF,
16'h175E, 16'hFFFF,
16'h175F, 16'hFFFF,
16'h1760, 16'hFFFF,
16'h1761, 16'hFFFF,
16'h1762, 16'hFFFF,
16'h1763, 16'hFFFF,
16'h1764, 16'hFFFF,
16'h1765, 16'hFFFF,
16'h1766, 16'hFFFF,
16'h1767, 16'hFFFF,
16'h1768, 16'hFFFF,
16'h1769, 16'hFFFF,
16'h176A, 16'hFFFF,
16'h176B, 16'hFFFF,
16'h176C, 16'hFFFF,
16'h176D, 16'hFFFF,
16'h176E, 16'hFFFF,
16'h176F, 16'hFFFF,
16'h1770, 16'hFFFF,
16'h1771, 16'hFFFF,
16'h1772, 16'hFFFF,
16'h1773, 16'hFFFF,
16'h1774, 16'hFFFF,
16'h1775, 16'hFFFF,
16'h1776, 16'hFFFF,
16'h1777, 16'hFFFF,
16'h1778, 16'hFFFF,
16'h1779, 16'hFFFF,
16'h177A, 16'hFFFF,
16'h177B, 16'hFFFF,
16'h177C, 16'hFFFF,
16'h177D, 16'hFFFF,
16'h177E, 16'hFFFF,
16'h177F, 16'hFFFF,
16'h1780, 16'hFFFF,
16'h1781, 16'hFFFF,
16'h1782, 16'hFFFF,
16'h1783, 16'hFFFF,
16'h1784, 16'hFFFF,
16'h1785, 16'hFFFF,
16'h1786, 16'hFFFF,
16'h1787, 16'hFFFF,
16'h1788, 16'hFFFF,
16'h1789, 16'hFFFF,
16'h178A, 16'hFFFF,
16'h178B, 16'hFFFF,
16'h178C, 16'hFFFF,
16'h178D, 16'hFFFF,
16'h178E, 16'hFFFF,
16'h178F, 16'hFFFF,
16'h1790, 16'hFFFF,
16'h1791, 16'hFFFF,
16'h1792, 16'hFFFF,
16'h1793, 16'hFFFF,
16'h1794, 16'hFFFF,
16'h1795, 16'hFFFF,
16'h1796, 16'hFFFF,
16'h1797, 16'hFFFF,
16'h1798, 16'hFFFF,
16'h1799, 16'hFFFF,
16'h179A, 16'hFFFF,
16'h179B, 16'hFFFF,
16'h179C, 16'hFFFF,
16'h179D, 16'hFFFF,
16'h179E, 16'hFFFF,
16'h179F, 16'hFFFF,
16'h17A0, 16'hFFFF,
16'h17A1, 16'hFFFF,
16'h17A2, 16'hFFFF,
16'h17A3, 16'hFFFF,
16'h17A4, 16'hFFFF,
16'h17A5, 16'hFFFF,
16'h17A6, 16'hFFFF,
16'h17A7, 16'hFFFF,
16'h17A8, 16'hFFFF,
16'h17A9, 16'hFFFF,
16'h17AA, 16'hFFFF,
16'h17AB, 16'hFFFF,
16'h17AC, 16'hFFFF,
16'h17AD, 16'hFFFF,
16'h17AE, 16'hFFFF,
16'h17AF, 16'hFFFF,
16'h17B0, 16'hFFFF,
16'h17B1, 16'hFFFF,
16'h17B2, 16'hFFFF,
16'h17B3, 16'hFFFF,
16'h17B4, 16'hFFFF,
16'h17B5, 16'hFFFF,
16'h17B6, 16'hFFFF,
16'h17B7, 16'hFFFF,
16'h17B8, 16'hFFFF,
16'h17B9, 16'hFFFF,
16'h17BA, 16'hFFFF,
16'h17BB, 16'hFFFF,
16'h17BC, 16'hFFFF,
16'h17BD, 16'hFFFF,
16'h17BE, 16'hFFFF,
16'h17BF, 16'hFFFF,
16'h17C0, 16'hFFFF,
16'h17C1, 16'hFFFF,
16'h17C2, 16'hFFFF,
16'h17C3, 16'hFFFF,
16'h17C4, 16'hFFFF,
16'h17C5, 16'hFFFF,
16'h17C6, 16'hFFFF,
16'h17C7, 16'hFFFF,
16'h17C8, 16'hFFFF,
16'h17C9, 16'hFFFF,
16'h17CA, 16'hFFFF,
16'h17CB, 16'hFFFF,
16'h17CC, 16'hFFFF,
16'h17CD, 16'hFFFF,
16'h17CE, 16'hFFFF,
16'h17CF, 16'hFFFF,
16'h17D0, 16'hFFFF,
16'h17D1, 16'hFFFF,
16'h17D2, 16'hFFFF,
16'h17D3, 16'hFFFF,
16'h17D4, 16'hFFFF,
16'h17D5, 16'hFFFF,
16'h17D6, 16'hFFFF,
16'h17D7, 16'hFFFF,
16'h17D8, 16'hFFFF,
16'h17D9, 16'hFFFF,
16'h17DA, 16'hFFFF,
16'h17DB, 16'hFFFF,
16'h17DC, 16'hFFFF,
16'h17DD, 16'hFFFF,
16'h17DE, 16'hFFFF,
16'h17DF, 16'hFFFF,
16'h17E0, 16'hFFFF,
16'h17E1, 16'hFFFF,
16'h17E2, 16'hFFFF,
16'h17E3, 16'hFFFF,
16'h17E4, 16'hFFFF,
16'h17E5, 16'hFFFF,
16'h17E6, 16'hFFFF,
16'h17E7, 16'hFFFF,
16'h17E8, 16'hFFFF,
16'h17E9, 16'hFFFF,
16'h17EA, 16'hFFFF,
16'h17EB, 16'hFFFF,
16'h17EC, 16'hFFFF,
16'h17ED, 16'hFFFF,
16'h17EE, 16'hFFFF,
16'h17EF, 16'hFFFF,
16'h17F0, 16'hFFFF,
16'h17F1, 16'hFFFF,
16'h17F2, 16'hFFFF,
16'h17F3, 16'hFFFF,
16'h17F4, 16'hFFFF,
16'h17F5, 16'hFFFF,
16'h17F6, 16'hFFFF,
16'h17F7, 16'hFFFF,
16'h17F8, 16'hFFFF,
16'h17F9, 16'hFFFF,
16'h17FA, 16'hFFFF,
16'h17FB, 16'hFFFF,
16'h17FC, 16'hFFFF,
16'h17FD, 16'hFFFF,
16'h17FE, 16'hFFFF,
16'h17FF, 16'hFFFF,
16'h1800, 16'hFFFF,
16'h1801, 16'hFFFF,
16'h1802, 16'hFFFF,
16'h1803, 16'hFFFF,
16'h1804, 16'hFFFF,
16'h1805, 16'hFFFF,
16'h1806, 16'hFFFF,
16'h1807, 16'hFFFF,
16'h1808, 16'hFFFF,
16'h1809, 16'hFFFF,
16'h180A, 16'hFFFF,
16'h180B, 16'hFFFF,
16'h180C, 16'hFFFF,
16'h180D, 16'hFFFF,
16'h180E, 16'hFFFF,
16'h180F, 16'hFFFF,
16'h1810, 16'hFFFF,
16'h1811, 16'hFFFF,
16'h1812, 16'hFFFF,
16'h1813, 16'hFFFF,
16'h1814, 16'hFFFF,
16'h1815, 16'hFFFF,
16'h1816, 16'hFFFF,
16'h1817, 16'hFFFF,
16'h1818, 16'hFFFF,
16'h1819, 16'hFFFF,
16'h181A, 16'hFFFF,
16'h181B, 16'hFFFF,
16'h181C, 16'hFFFF,
16'h181D, 16'hFFFF,
16'h181E, 16'hFFFF,
16'h181F, 16'hFFFF,
16'h1820, 16'hFFFF,
16'h1821, 16'hFFFF,
16'h1822, 16'hFFFF,
16'h1823, 16'hFFFF,
16'h1824, 16'hFFFF,
16'h1825, 16'hFFFF,
16'h1826, 16'hFFFF,
16'h1827, 16'hFFFF,
16'h1828, 16'hFFFF,
16'h1829, 16'hFFFF,
16'h182A, 16'hFFFF,
16'h182B, 16'hFFFF,
16'h182C, 16'hFFFF,
16'h182D, 16'hFFFF,
16'h182E, 16'hFFFF,
16'h182F, 16'hFFFF,
16'h1830, 16'hFFFF,
16'h1831, 16'hFFFF,
16'h1832, 16'hFFFF,
16'h1833, 16'hFFFF,
16'h1834, 16'hFFFF,
16'h1835, 16'hFFFF,
16'h1836, 16'hFFFF,
16'h1837, 16'hFFFF,
16'h1838, 16'hFFFF,
16'h1839, 16'hFFFF,
16'h183A, 16'hFFFF,
16'h183B, 16'hFFFF,
16'h183C, 16'hFFFF,
16'h183D, 16'hFFFF,
16'h183E, 16'hFFFF,
16'h183F, 16'hFFFF,
16'h1840, 16'hFFFF,
16'h1841, 16'hFFFF,
16'h1842, 16'hFFFF,
16'h1843, 16'hFFFF,
16'h1844, 16'hFFFF,
16'h1845, 16'hFFFF,
16'h1846, 16'hFFFF,
16'h1847, 16'hFFFF,
16'h1848, 16'hFFFF,
16'h1849, 16'hFFFF,
16'h184A, 16'hFFFF,
16'h184B, 16'hFFFF,
16'h184C, 16'hFFFF,
16'h184D, 16'hFFFF,
16'h184E, 16'hFFFF,
16'h184F, 16'hFFFF,
16'h1850, 16'hFFFF,
16'h1851, 16'hFFFF,
16'h1852, 16'hFFFF,
16'h1853, 16'hFFFF,
16'h1854, 16'hFFFF,
16'h1855, 16'hFFFF,
16'h1856, 16'hFFFF,
16'h1857, 16'hFFFF,
16'h1858, 16'hFFFF,
16'h1859, 16'hFFFF,
16'h185A, 16'hFFFF,
16'h185B, 16'hFFFF,
16'h185C, 16'hFFFF,
16'h185D, 16'hFFFF,
16'h185E, 16'hFFFF,
16'h185F, 16'hFFFF,
16'h1860, 16'hFFFF,
16'h1861, 16'hFFFF,
16'h1862, 16'hFFFF,
16'h1863, 16'hFFFF,
16'h1864, 16'hFFFF,
16'h1865, 16'hFFFF,
16'h1866, 16'hFFFF,
16'h1867, 16'hFFFF,
16'h1868, 16'hFFFF,
16'h1869, 16'hFFFF,
16'h186A, 16'hFFFF,
16'h186B, 16'hFFFF,
16'h186C, 16'hFFFF,
16'h186D, 16'hFFFF,
16'h186E, 16'hFFFF,
16'h186F, 16'hFFFF,
16'h1870, 16'hFFFF,
16'h1871, 16'hFFFF,
16'h1872, 16'hFFFF,
16'h1873, 16'hFFFF,
16'h1874, 16'hFFFF,
16'h1875, 16'hFFFF,
16'h1876, 16'hFFFF,
16'h1877, 16'hFFFF,
16'h1878, 16'hFFFF,
16'h1879, 16'hFFFF,
16'h187A, 16'hFFFF,
16'h187B, 16'hFFFF,
16'h187C, 16'hFFFF,
16'h187D, 16'hFFFF,
16'h187E, 16'hFFFF,
16'h187F, 16'hFFFF,
16'h1880, 16'hFFFF,
16'h1881, 16'hFFFF,
16'h1882, 16'hFFFF,
16'h1883, 16'hFFFF,
16'h1884, 16'hFFFF,
16'h1885, 16'hFFFF,
16'h1886, 16'hFFFF,
16'h1887, 16'hFFFF,
16'h1888, 16'hFFFF,
16'h1889, 16'hFFFF,
16'h188A, 16'hFFFF,
16'h188B, 16'hFFFF,
16'h188C, 16'hFFFF,
16'h188D, 16'hFFFF,
16'h188E, 16'hFFFF,
16'h188F, 16'hFFFF,
16'h1890, 16'hFFFF,
16'h1891, 16'hFFFF,
16'h1892, 16'hFFFF,
16'h1893, 16'hFFFF,
16'h1894, 16'hFFFF,
16'h1895, 16'hFFFF,
16'h1896, 16'hFFFF,
16'h1897, 16'hFFFF,
16'h1898, 16'hFFFF,
16'h1899, 16'hFFFF,
16'h189A, 16'hFFFF,
16'h189B, 16'hFFFF,
16'h189C, 16'hFFFF,
16'h189D, 16'hFFFF,
16'h189E, 16'hFFFF,
16'h189F, 16'hFFFF,
16'h18A0, 16'hFFFF,
16'h18A1, 16'hFFFF,
16'h18A2, 16'hFFFF,
16'h18A3, 16'hFFFF,
16'h18A4, 16'hFFFF,
16'h18A5, 16'hFFFF,
16'h18A6, 16'hFFFF,
16'h18A7, 16'hFFFF,
16'h18A8, 16'hFFFF,
16'h18A9, 16'hFFFF,
16'h18AA, 16'hFFFF,
16'h18AB, 16'hFFFF,
16'h18AC, 16'hFFFF,
16'h18AD, 16'hFFFF,
16'h18AE, 16'hFFFF,
16'h18AF, 16'hFFFF,
16'h18B0, 16'hFFFF,
16'h18B1, 16'hFFFF,
16'h18B2, 16'hFFFF,
16'h18B3, 16'hFFFF,
16'h18B4, 16'hFFFF,
16'h18B5, 16'hFFFF,
16'h18B6, 16'hFFFF,
16'h18B7, 16'hFFFF,
16'h18B8, 16'hFFFF,
16'h18B9, 16'hFFFF,
16'h18BA, 16'hFFFF,
16'h18BB, 16'hFFFF,
16'h18BC, 16'hFFFF,
16'h18BD, 16'hFFFF,
16'h18BE, 16'hFFFF,
16'h18BF, 16'hFFFF,
16'h18C0, 16'hFFFF,
16'h18C1, 16'hFFFF,
16'h18C2, 16'hFFFF,
16'h18C3, 16'hFFFF,
16'h18C4, 16'hFFFF,
16'h18C5, 16'hFFFF,
16'h18C6, 16'hFFFF,
16'h18C7, 16'hFFFF,
16'h18C8, 16'hFFFF,
16'h18C9, 16'hFFFF,
16'h18CA, 16'hFFFF,
16'h18CB, 16'hFFFF,
16'h18CC, 16'hFFFF,
16'h18CD, 16'hFFFF,
16'h18CE, 16'hFFFF,
16'h18CF, 16'hFFFF,
16'h18D0, 16'hFFFF,
16'h18D1, 16'hFFFF,
16'h18D2, 16'hFFFF,
16'h18D3, 16'hFFFF,
16'h18D4, 16'hFFFF,
16'h18D5, 16'hFFFF,
16'h18D6, 16'hFFFF,
16'h18D7, 16'hFFFF,
16'h18D8, 16'hFFFF,
16'h18D9, 16'hFFFF,
16'h18DA, 16'hFFFF,
16'h18DB, 16'hFFFF,
16'h18DC, 16'hFFFF,
16'h18DD, 16'hFFFF,
16'h18DE, 16'hFFFF,
16'h18DF, 16'hFFFF,
16'h18E0, 16'hFFFF,
16'h18E1, 16'hFFFF,
16'h18E2, 16'hFFFF,
16'h18E3, 16'hFFFF,
16'h18E4, 16'hFFFF,
16'h18E5, 16'hFFFF,
16'h18E6, 16'hFFFF,
16'h18E7, 16'hFFFF,
16'h18E8, 16'hFFFF,
16'h18E9, 16'hFFFF,
16'h18EA, 16'hFFFF,
16'h18EB, 16'hFFFF,
16'h18EC, 16'hFFFF,
16'h18ED, 16'hFFFF,
16'h18EE, 16'hFFFF,
16'h18EF, 16'hFFFF,
16'h18F0, 16'hFFFF,
16'h18F1, 16'hFFFF,
16'h18F2, 16'hFFFF,
16'h18F3, 16'hFFFF,
16'h18F4, 16'hFFFF,
16'h18F5, 16'hFFFF,
16'h18F6, 16'hFFFF,
16'h18F7, 16'hFFFF,
16'h18F8, 16'hFFFF,
16'h18F9, 16'hFFFF,
16'h18FA, 16'hFFFF,
16'h18FB, 16'hFFFF,
16'h18FC, 16'hFFFF,
16'h18FD, 16'hFFFF,
16'h18FE, 16'hFFFF,
16'h18FF, 16'hFFFF,
16'h1900, 16'hFFFF,
16'h1901, 16'hFFFF,
16'h1902, 16'hFFFF,
16'h1903, 16'hFFFF,
16'h1904, 16'hFFFF,
16'h1905, 16'hFFFF,
16'h1906, 16'hFFFF,
16'h1907, 16'hFFFF,
16'h1908, 16'hFFFF,
16'h1909, 16'hFFFF,
16'h190A, 16'hFFFF,
16'h190B, 16'hFFFF,
16'h190C, 16'hFFFF,
16'h190D, 16'hFFFF,
16'h190E, 16'hFFFF,
16'h190F, 16'hFFFF,
16'h1910, 16'hFFFF,
16'h1911, 16'hFFFF,
16'h1912, 16'hFFFF,
16'h1913, 16'hFFFF,
16'h1914, 16'hFFFF,
16'h1915, 16'hFFFF,
16'h1916, 16'hFFFF,
16'h1917, 16'hFFFF,
16'h1918, 16'hFFFF,
16'h1919, 16'hFFFF,
16'h191A, 16'hFFFF,
16'h191B, 16'hFFFF,
16'h191C, 16'hFFFF,
16'h191D, 16'hFFFF,
16'h191E, 16'hFFFF,
16'h191F, 16'hFFFF,
16'h1920, 16'hFFFF,
16'h1921, 16'hFFFF,
16'h1922, 16'hFFFF,
16'h1923, 16'hFFFF,
16'h1924, 16'hFFFF,
16'h1925, 16'hFFFF,
16'h1926, 16'hFFFF,
16'h1927, 16'hFFFF,
16'h1928, 16'hFFFF,
16'h1929, 16'hFFFF,
16'h192A, 16'hFFFF,
16'h192B, 16'hFFFF,
16'h192C, 16'hFFFF,
16'h192D, 16'hFFFF,
16'h192E, 16'hFFFF,
16'h192F, 16'hFFFF,
16'h1930, 16'hFFFF,
16'h1931, 16'hFFFF,
16'h1932, 16'hFFFF,
16'h1933, 16'hFFFF,
16'h1934, 16'hFFFF,
16'h1935, 16'hFFFF,
16'h1936, 16'hFFFF,
16'h1937, 16'hFFFF,
16'h1938, 16'hFFFF,
16'h1939, 16'hFFFF,
16'h193A, 16'hFFFF,
16'h193B, 16'hFFFF,
16'h193C, 16'hFFFF,
16'h193D, 16'hFFFF,
16'h193E, 16'hFFFF,
16'h193F, 16'hFFFF,
16'h1940, 16'hFFFF,
16'h1941, 16'hFFFF,
16'h1942, 16'hFFFF,
16'h1943, 16'hFFFF,
16'h1944, 16'hFFFF,
16'h1945, 16'hFFFF,
16'h1946, 16'hFFFF,
16'h1947, 16'hFFFF,
16'h1948, 16'hFFFF,
16'h1949, 16'hFFFF,
16'h194A, 16'hFFFF,
16'h194B, 16'hFFFF,
16'h194C, 16'hFFFF,
16'h194D, 16'hFFFF,
16'h194E, 16'hFFFF,
16'h194F, 16'hFFFF,
16'h1950, 16'hFFFF,
16'h1951, 16'hFFFF,
16'h1952, 16'hFFFF,
16'h1953, 16'hFFFF,
16'h1954, 16'hFFFF,
16'h1955, 16'hFFFF,
16'h1956, 16'hFFFF,
16'h1957, 16'hFFFF,
16'h1958, 16'hFFFF,
16'h1959, 16'hFFFF,
16'h195A, 16'hFFFF,
16'h195B, 16'hFFFF,
16'h195C, 16'hFFFF,
16'h195D, 16'hFFFF,
16'h195E, 16'hFFFF,
16'h195F, 16'hFFFF,
16'h1960, 16'hFFFF,
16'h1961, 16'hFFFF,
16'h1962, 16'hFFFF,
16'h1963, 16'hFFFF,
16'h1964, 16'hFFFF,
16'h1965, 16'hFFFF,
16'h1966, 16'hFFFF,
16'h1967, 16'hFFFF,
16'h1968, 16'hFFFF,
16'h1969, 16'hFFFF,
16'h196A, 16'hFFFF,
16'h196B, 16'hFFFF,
16'h196C, 16'hFFFF,
16'h196D, 16'hFFFF,
16'h196E, 16'hFFFF,
16'h196F, 16'hFFFF,
16'h1970, 16'hFFFF,
16'h1971, 16'hFFFF,
16'h1972, 16'hFFFF,
16'h1973, 16'hFFFF,
16'h1974, 16'hFFFF,
16'h1975, 16'hFFFF,
16'h1976, 16'hFFFF,
16'h1977, 16'hFFFF,
16'h1978, 16'hFFFF,
16'h1979, 16'hFFFF,
16'h197A, 16'hFFFF,
16'h197B, 16'hFFFF,
16'h197C, 16'hFFFF,
16'h197D, 16'hFFFF,
16'h197E, 16'hFFFF,
16'h197F, 16'hFFFF,
16'h1980, 16'hFFFF,
16'h1981, 16'hFFFF,
16'h1982, 16'hFFFF,
16'h1983, 16'hFFFF,
16'h1984, 16'hFFFF,
16'h1985, 16'hFFFF,
16'h1986, 16'hFFFF,
16'h1987, 16'hFFFF,
16'h1988, 16'hFFFF,
16'h1989, 16'hFFFF,
16'h198A, 16'hFFFF,
16'h198B, 16'hFFFF,
16'h198C, 16'hFFFF,
16'h198D, 16'hFFFF,
16'h198E, 16'hFFFF,
16'h198F, 16'hFFFF,
16'h1990, 16'hFFFF,
16'h1991, 16'hFFFF,
16'h1992, 16'hFFFF,
16'h1993, 16'hFFFF,
16'h1994, 16'hFFFF,
16'h1995, 16'hFFFF,
16'h1996, 16'hFFFF,
16'h1997, 16'hFFFF,
16'h1998, 16'hFFFF,
16'h1999, 16'hFFFF,
16'h199A, 16'hFFFF,
16'h199B, 16'hFFFF,
16'h199C, 16'hFFFF,
16'h199D, 16'hFFFF,
16'h199E, 16'hFFFF,
16'h199F, 16'hFFFF,
16'h19A0, 16'hFFFF,
16'h19A1, 16'hFFFF,
16'h19A2, 16'hFFFF,
16'h19A3, 16'hFFFF,
16'h19A4, 16'hFFFF,
16'h19A5, 16'hFFFF,
16'h19A6, 16'hFFFF,
16'h19A7, 16'hFFFF,
16'h19A8, 16'hFFFF,
16'h19A9, 16'hFFFF,
16'h19AA, 16'hFFFF,
16'h19AB, 16'hFFFF,
16'h19AC, 16'hFFFF,
16'h19AD, 16'hFFFF,
16'h19AE, 16'hFFFF,
16'h19AF, 16'hFFFF,
16'h19B0, 16'hFFFF,
16'h19B1, 16'hFFFF,
16'h19B2, 16'hFFFF,
16'h19B3, 16'hFFFF,
16'h19B4, 16'hFFFF,
16'h19B5, 16'hFFFF,
16'h19B6, 16'hFFFF,
16'h19B7, 16'hFFFF,
16'h19B8, 16'hFFFF,
16'h19B9, 16'hFFFF,
16'h19BA, 16'hFFFF,
16'h19BB, 16'hFFFF,
16'h19BC, 16'hFFFF,
16'h19BD, 16'hFFFF,
16'h19BE, 16'hFFFF,
16'h19BF, 16'hFFFF,
16'h19C0, 16'hFFFF,
16'h19C1, 16'hFFFF,
16'h19C2, 16'hFFFF,
16'h19C3, 16'hFFFF,
16'h19C4, 16'hFFFF,
16'h19C5, 16'hFFFF,
16'h19C6, 16'hFFFF,
16'h19C7, 16'hFFFF,
16'h19C8, 16'hFFFF,
16'h19C9, 16'hFFFF,
16'h19CA, 16'hFFFF,
16'h19CB, 16'hFFFF,
16'h19CC, 16'hFFFF,
16'h19CD, 16'hFFFF,
16'h19CE, 16'hFFFF,
16'h19CF, 16'hFFFF,
16'h19D0, 16'hFFFF,
16'h19D1, 16'hFFFF,
16'h19D2, 16'hFFFF,
16'h19D3, 16'hFFFF,
16'h19D4, 16'hFFFF,
16'h19D5, 16'hFFFF,
16'h19D6, 16'hFFFF,
16'h19D7, 16'hFFFF,
16'h19D8, 16'hFFFF,
16'h19D9, 16'hFFFF,
16'h19DA, 16'hFFFF,
16'h19DB, 16'hFFFF,
16'h19DC, 16'hFFFF,
16'h19DD, 16'hFFFF,
16'h19DE, 16'hFFFF,
16'h19DF, 16'hFFFF,
16'h19E0, 16'hFFFF,
16'h19E1, 16'hFFFF,
16'h19E2, 16'hFFFF,
16'h19E3, 16'hFFFF,
16'h19E4, 16'hFFFF,
16'h19E5, 16'hFFFF,
16'h19E6, 16'hFFFF,
16'h19E7, 16'hFFFF,
16'h19E8, 16'hFFFF,
16'h19E9, 16'hFFFF,
16'h19EA, 16'hFFFF,
16'h19EB, 16'hFFFF,
16'h19EC, 16'hFFFF,
16'h19ED, 16'hFFFF,
16'h19EE, 16'hFFFF,
16'h19EF, 16'hFFFF,
16'h19F0, 16'hFFFF,
16'h19F1, 16'hFFFF,
16'h19F2, 16'hFFFF,
16'h19F3, 16'hFFFF,
16'h19F4, 16'hFFFF,
16'h19F5, 16'hFFFF,
16'h19F6, 16'hFFFF,
16'h19F7, 16'hFFFF,
16'h19F8, 16'hFFFF,
16'h19F9, 16'hFFFF,
16'h19FA, 16'hFFFF,
16'h19FB, 16'hFFFF,
16'h19FC, 16'hFFFF,
16'h19FD, 16'hFFFF,
16'h19FE, 16'hFFFF,
16'h19FF, 16'hFFFF,
16'h1A00, 16'hFFFF,
16'h1A01, 16'hFFFF,
16'h1A02, 16'hFFFF,
16'h1A03, 16'hFFFF,
16'h1A04, 16'hFFFF,
16'h1A05, 16'hFFFF,
16'h1A06, 16'hFFFF,
16'h1A07, 16'hFFFF,
16'h1A08, 16'hFFFF,
16'h1A09, 16'hFFFF,
16'h1A0A, 16'hFFFF,
16'h1A0B, 16'hFFFF,
16'h1A0C, 16'hFFFF,
16'h1A0D, 16'hFFFF,
16'h1A0E, 16'hFFFF,
16'h1A0F, 16'hFFFF,
16'h1A10, 16'hFFFF,
16'h1A11, 16'hFFFF,
16'h1A12, 16'hFFFF,
16'h1A13, 16'hFFFF,
16'h1A14, 16'hFFFF,
16'h1A15, 16'hFFFF,
16'h1A16, 16'hFFFF,
16'h1A17, 16'hFFFF,
16'h1A18, 16'hFFFF,
16'h1A19, 16'hFFFF,
16'h1A1A, 16'hFFFF,
16'h1A1B, 16'hFFFF,
16'h1A1C, 16'hFFFF,
16'h1A1D, 16'hFFFF,
16'h1A1E, 16'hFFFF,
16'h1A1F, 16'hFFFF,
16'h1A20, 16'hFFFF,
16'h1A21, 16'hFFFF,
16'h1A22, 16'hFFFF,
16'h1A23, 16'hFFFF,
16'h1A24, 16'hFFFF,
16'h1A25, 16'hFFFF,
16'h1A26, 16'hFFFF,
16'h1A27, 16'hFFFF,
16'h1A28, 16'hFFFF,
16'h1A29, 16'hFFFF,
16'h1A2A, 16'hFFFF,
16'h1A2B, 16'hFFFF,
16'h1A2C, 16'hFFFF,
16'h1A2D, 16'hFFFF,
16'h1A2E, 16'hFFFF,
16'h1A2F, 16'hFFFF,
16'h1A30, 16'hFFFF,
16'h1A31, 16'hFFFF,
16'h1A32, 16'hFFFF,
16'h1A33, 16'hFFFF,
16'h1A34, 16'hFFFF,
16'h1A35, 16'hFFFF,
16'h1A36, 16'hFFFF,
16'h1A37, 16'hFFFF,
16'h1A38, 16'hFFFF,
16'h1A39, 16'hFFFF,
16'h1A3A, 16'hFFFF,
16'h1A3B, 16'hFFFF,
16'h1A3C, 16'hFFFF,
16'h1A3D, 16'hFFFF,
16'h1A3E, 16'hFFFF,
16'h1A3F, 16'hFFFF,
16'h1A40, 16'hFFFF,
16'h1A41, 16'hFFFF,
16'h1A42, 16'hFFFF,
16'h1A43, 16'hFFFF,
16'h1A44, 16'hFFFF,
16'h1A45, 16'hFFFF,
16'h1A46, 16'hFFFF,
16'h1A47, 16'hFFFF,
16'h1A48, 16'hFFFF,
16'h1A49, 16'hFFFF,
16'h1A4A, 16'hFFFF,
16'h1A4B, 16'hFFFF,
16'h1A4C, 16'hFFFF,
16'h1A4D, 16'hFFFF,
16'h1A4E, 16'hFFFF,
16'h1A4F, 16'hFFFF,
16'h1A50, 16'hFFFF,
16'h1A51, 16'hFFFF,
16'h1A52, 16'hFFFF,
16'h1A53, 16'hFFFF,
16'h1A54, 16'hFFFF,
16'h1A55, 16'hFFFF,
16'h1A56, 16'hFFFF,
16'h1A57, 16'hFFFF,
16'h1A58, 16'hFFFF,
16'h1A59, 16'hFFFF,
16'h1A5A, 16'hFFFF,
16'h1A5B, 16'hFFFF,
16'h1A5C, 16'hFFFF,
16'h1A5D, 16'hFFFF,
16'h1A5E, 16'hFFFF,
16'h1A5F, 16'hFFFF,
16'h1A60, 16'hFFFF,
16'h1A61, 16'hFFFF,
16'h1A62, 16'hFFFF,
16'h1A63, 16'hFFFF,
16'h1A64, 16'hFFFF,
16'h1A65, 16'hFFFF,
16'h1A66, 16'hFFFF,
16'h1A67, 16'hFFFF,
16'h1A68, 16'hFFFF,
16'h1A69, 16'hFFFF,
16'h1A6A, 16'hFFFF,
16'h1A6B, 16'hFFFF,
16'h1A6C, 16'hFFFF,
16'h1A6D, 16'hFFFF,
16'h1A6E, 16'hFFFF,
16'h1A6F, 16'hFFFF,
16'h1A70, 16'hFFFF,
16'h1A71, 16'hFFFF,
16'h1A72, 16'hFFFF,
16'h1A73, 16'hFFFF,
16'h1A74, 16'hFFFF,
16'h1A75, 16'hFFFF,
16'h1A76, 16'hFFFF,
16'h1A77, 16'hFFFF,
16'h1A78, 16'hFFFF,
16'h1A79, 16'hFFFF,
16'h1A7A, 16'hFFFF,
16'h1A7B, 16'hFFFF,
16'h1A7C, 16'hFFFF,
16'h1A7D, 16'hFFFF,
16'h1A7E, 16'hFFFF,
16'h1A7F, 16'hFFFF,
16'h1A80, 16'hFFFF,
16'h1A81, 16'hFFFF,
16'h1A82, 16'hFFFF,
16'h1A83, 16'hFFFF,
16'h1A84, 16'hFFFF,
16'h1A85, 16'hFFFF,
16'h1A86, 16'hFFFF,
16'h1A87, 16'hFFFF,
16'h1A88, 16'hFFFF,
16'h1A89, 16'hFFFF,
16'h1A8A, 16'hFFFF,
16'h1A8B, 16'hFFFF,
16'h1A8C, 16'hFFFF,
16'h1A8D, 16'hFFFF,
16'h1A8E, 16'hFFFF,
16'h1A8F, 16'hFFFF,
16'h1A90, 16'hFFFF,
16'h1A91, 16'hFFFF,
16'h1A92, 16'hFFFF,
16'h1A93, 16'hFFFF,
16'h1A94, 16'hFFFF,
16'h1A95, 16'hFFFF,
16'h1A96, 16'hFFFF,
16'h1A97, 16'hFFFF,
16'h1A98, 16'hFFFF,
16'h1A99, 16'hFFFF,
16'h1A9A, 16'hFFFF,
16'h1A9B, 16'hFFFF,
16'h1A9C, 16'hFFFF,
16'h1A9D, 16'hFFFF,
16'h1A9E, 16'hFFFF,
16'h1A9F, 16'hFFFF,
16'h1AA0, 16'hFFFF,
16'h1AA1, 16'hFFFF,
16'h1AA2, 16'hFFFF,
16'h1AA3, 16'hFFFF,
16'h1AA4, 16'hFFFF,
16'h1AA5, 16'hFFFF,
16'h1AA6, 16'hFFFF,
16'h1AA7, 16'hFFFF,
16'h1AA8, 16'hFFFF,
16'h1AA9, 16'hFFFF,
16'h1AAA, 16'hFFFF,
16'h1AAB, 16'hFFFF,
16'h1AAC, 16'hFFFF,
16'h1AAD, 16'hFFFF,
16'h1AAE, 16'hFFFF,
16'h1AAF, 16'hFFFF,
16'h1AB0, 16'hFFFF,
16'h1AB1, 16'hFFFF,
16'h1AB2, 16'hFFFF,
16'h1AB3, 16'hFFFF,
16'h1AB4, 16'hFFFF,
16'h1AB5, 16'hFFFF,
16'h1AB6, 16'hFFFF,
16'h1AB7, 16'hFFFF,
16'h1AB8, 16'hFFFF,
16'h1AB9, 16'hFFFF,
16'h1ABA, 16'hFFFF,
16'h1ABB, 16'hFFFF,
16'h1ABC, 16'hFFFF,
16'h1ABD, 16'hFFFF,
16'h1ABE, 16'hFFFF,
16'h1ABF, 16'hFFFF,
16'h1AC0, 16'hFFFF,
16'h1AC1, 16'hFFFF,
16'h1AC2, 16'hFFFF,
16'h1AC3, 16'hFFFF,
16'h1AC4, 16'hFFFF,
16'h1AC5, 16'hFFFF,
16'h1AC6, 16'hFFFF,
16'h1AC7, 16'hFFFF,
16'h1AC8, 16'hFFFF,
16'h1AC9, 16'hFFFF,
16'h1ACA, 16'hFFFF,
16'h1ACB, 16'hFFFF,
16'h1ACC, 16'hFFFF,
16'h1ACD, 16'hFFFF,
16'h1ACE, 16'hFFFF,
16'h1ACF, 16'hFFFF,
16'h1AD0, 16'hFFFF,
16'h1AD1, 16'hFFFF,
16'h1AD2, 16'hFFFF,
16'h1AD3, 16'hFFFF,
16'h1AD4, 16'hFFFF,
16'h1AD5, 16'hFFFF,
16'h1AD6, 16'hFFFF,
16'h1AD7, 16'hFFFF,
16'h1AD8, 16'hFFFF,
16'h1AD9, 16'hFFFF,
16'h1ADA, 16'hFFFF,
16'h1ADB, 16'hFFFF,
16'h1ADC, 16'hFFFF,
16'h1ADD, 16'hFFFF,
16'h1ADE, 16'hFFFF,
16'h1ADF, 16'hFFFF,
16'h1AE0, 16'hFFFF,
16'h1AE1, 16'hFFFF,
16'h1AE2, 16'hFFFF,
16'h1AE3, 16'hFFFF,
16'h1AE4, 16'hFFFF,
16'h1AE5, 16'hFFFF,
16'h1AE6, 16'hFFFF,
16'h1AE7, 16'hFFFF,
16'h1AE8, 16'hFFFF,
16'h1AE9, 16'hFFFF,
16'h1AEA, 16'hFFFF,
16'h1AEB, 16'hFFFF,
16'h1AEC, 16'hFFFF,
16'h1AED, 16'hFFFF,
16'h1AEE, 16'hFFFF,
16'h1AEF, 16'hFFFF,
16'h1AF0, 16'hFFFF,
16'h1AF1, 16'hFFFF,
16'h1AF2, 16'hFFFF,
16'h1AF3, 16'hFFFF,
16'h1AF4, 16'hFFFF,
16'h1AF5, 16'hFFFF,
16'h1AF6, 16'hFFFF,
16'h1AF7, 16'hFFFF,
16'h1AF8, 16'hFFFF,
16'h1AF9, 16'hFFFF,
16'h1AFA, 16'hFFFF,
16'h1AFB, 16'hFFFF,
16'h1AFC, 16'hFFFF,
16'h1AFD, 16'hFFFF,
16'h1AFE, 16'hFFFF,
16'h1AFF, 16'hFFFF,
16'h1B00, 16'hFFFF,
16'h1B01, 16'hFFFF,
16'h1B02, 16'hFFFF,
16'h1B03, 16'hFFFF,
16'h1B04, 16'hFFFF,
16'h1B05, 16'hFFFF,
16'h1B06, 16'hFFFF,
16'h1B07, 16'hFFFF,
16'h1B08, 16'hFFFF,
16'h1B09, 16'hFFFF,
16'h1B0A, 16'hFFFF,
16'h1B0B, 16'hFFFF,
16'h1B0C, 16'hFFFF,
16'h1B0D, 16'hFFFF,
16'h1B0E, 16'hFFFF,
16'h1B0F, 16'hFFFF,
16'h1B10, 16'hFFFF,
16'h1B11, 16'hFFFF,
16'h1B12, 16'hFFFF,
16'h1B13, 16'hFFFF,
16'h1B14, 16'hFFFF,
16'h1B15, 16'hFFFF,
16'h1B16, 16'hFFFF,
16'h1B17, 16'hFFFF,
16'h1B18, 16'hFFFF,
16'h1B19, 16'hFFFF,
16'h1B1A, 16'hFFFF,
16'h1B1B, 16'hFFFF,
16'h1B1C, 16'hFFFF,
16'h1B1D, 16'hFFFF,
16'h1B1E, 16'hFFFF,
16'h1B1F, 16'hFFFF,
16'h1B20, 16'hFFFF,
16'h1B21, 16'hFFFF,
16'h1B22, 16'hFFFF,
16'h1B23, 16'hFFFF,
16'h1B24, 16'hFFFF,
16'h1B25, 16'hFFFF,
16'h1B26, 16'hFFFF,
16'h1B27, 16'hFFFF,
16'h1B28, 16'hFFFF,
16'h1B29, 16'hFFFF,
16'h1B2A, 16'hFFFF,
16'h1B2B, 16'hFFFF,
16'h1B2C, 16'hFFFF,
16'h1B2D, 16'hFFFF,
16'h1B2E, 16'hFFFF,
16'h1B2F, 16'hFFFF,
16'h1B30, 16'hFFFF,
16'h1B31, 16'hFFFF,
16'h1B32, 16'hFFFF,
16'h1B33, 16'hFFFF,
16'h1B34, 16'hFFFF,
16'h1B35, 16'hFFFF,
16'h1B36, 16'hFFFF,
16'h1B37, 16'hFFFF,
16'h1B38, 16'hFFFF,
16'h1B39, 16'hFFFF,
16'h1B3A, 16'hFFFF,
16'h1B3B, 16'hFFFF,
16'h1B3C, 16'hFFFF,
16'h1B3D, 16'hFFFF,
16'h1B3E, 16'hFFFF,
16'h1B3F, 16'hFFFF,
16'h1B40, 16'hFFFF,
16'h1B41, 16'hFFFF,
16'h1B42, 16'hFFFF,
16'h1B43, 16'hFFFF,
16'h1B44, 16'hFFFF,
16'h1B45, 16'hFFFF,
16'h1B46, 16'hFFFF,
16'h1B47, 16'hFFFF,
16'h1B48, 16'hFFFF,
16'h1B49, 16'hFFFF,
16'h1B4A, 16'hFFFF,
16'h1B4B, 16'hFFFF,
16'h1B4C, 16'hFFFF,
16'h1B4D, 16'hFFFF,
16'h1B4E, 16'hFFFF,
16'h1B4F, 16'hFFFF,
16'h1B50, 16'hFFFF,
16'h1B51, 16'hFFFF,
16'h1B52, 16'hFFFF,
16'h1B53, 16'hFFFF,
16'h1B54, 16'hFFFF,
16'h1B55, 16'hFFFF,
16'h1B56, 16'hFFFF,
16'h1B57, 16'hFFFF,
16'h1B58, 16'hFFFF,
16'h1B59, 16'hFFFF,
16'h1B5A, 16'hFFFF,
16'h1B5B, 16'hFFFF,
16'h1B5C, 16'hFFFF,
16'h1B5D, 16'hFFFF,
16'h1B5E, 16'hFFFF,
16'h1B5F, 16'hFFFF,
16'h1B60, 16'hFFFF,
16'h1B61, 16'hFFFF,
16'h1B62, 16'hFFFF,
16'h1B63, 16'hFFFF,
16'h1B64, 16'hFFFF,
16'h1B65, 16'hFFFF,
16'h1B66, 16'hFFFF,
16'h1B67, 16'hFFFF,
16'h1B68, 16'hFFFF,
16'h1B69, 16'hFFFF,
16'h1B6A, 16'hFFFF,
16'h1B6B, 16'hFFFF,
16'h1B6C, 16'hFFFF,
16'h1B6D, 16'hFFFF,
16'h1B6E, 16'hFFFF,
16'h1B6F, 16'hFFFF,
16'h1B70, 16'hFFFF,
16'h1B71, 16'hFFFF,
16'h1B72, 16'hFFFF,
16'h1B73, 16'hFFFF,
16'h1B74, 16'hFFFF,
16'h1B75, 16'hFFFF,
16'h1B76, 16'hFFFF,
16'h1B77, 16'hFFFF,
16'h1B78, 16'hFFFF,
16'h1B79, 16'hFFFF,
16'h1B7A, 16'hFFFF,
16'h1B7B, 16'hFFFF,
16'h1B7C, 16'hFFFF,
16'h1B7D, 16'hFFFF,
16'h1B7E, 16'hFFFF,
16'h1B7F, 16'hFFFF,
16'h1B80, 16'hFFFF,
16'h1B81, 16'hFFFF,
16'h1B82, 16'hFFFF,
16'h1B83, 16'hFFFF,
16'h1B84, 16'hFFFF,
16'h1B85, 16'hFFFF,
16'h1B86, 16'hFFFF,
16'h1B87, 16'hFFFF,
16'h1B88, 16'hFFFF,
16'h1B89, 16'hFFFF,
16'h1B8A, 16'hFFFF,
16'h1B8B, 16'hFFFF,
16'h1B8C, 16'hFFFF,
16'h1B8D, 16'hFFFF,
16'h1B8E, 16'hFFFF,
16'h1B8F, 16'hFFFF,
16'h1B90, 16'hFFFF,
16'h1B91, 16'hFFFF,
16'h1B92, 16'hFFFF,
16'h1B93, 16'hFFFF,
16'h1B94, 16'hFFFF,
16'h1B95, 16'hFFFF,
16'h1B96, 16'hFFFF,
16'h1B97, 16'hFFFF,
16'h1B98, 16'hFFFF,
16'h1B99, 16'hFFFF,
16'h1B9A, 16'hFFFF,
16'h1B9B, 16'hFFFF,
16'h1B9C, 16'hFFFF,
16'h1B9D, 16'hFFFF,
16'h1B9E, 16'hFFFF,
16'h1B9F, 16'hFFFF,
16'h1BA0, 16'hFFFF,
16'h1BA1, 16'hFFFF,
16'h1BA2, 16'hFFFF,
16'h1BA3, 16'hFFFF,
16'h1BA4, 16'hFFFF,
16'h1BA5, 16'hFFFF,
16'h1BA6, 16'hFFFF,
16'h1BA7, 16'hFFFF,
16'h1BA8, 16'hFFFF,
16'h1BA9, 16'hFFFF,
16'h1BAA, 16'hFFFF,
16'h1BAB, 16'hFFFF,
16'h1BAC, 16'hFFFF,
16'h1BAD, 16'hFFFF,
16'h1BAE, 16'hFFFF,
16'h1BAF, 16'hFFFF,
16'h1BB0, 16'hFFFF,
16'h1BB1, 16'hFFFF,
16'h1BB2, 16'hFFFF,
16'h1BB3, 16'hFFFF,
16'h1BB4, 16'hFFFF,
16'h1BB5, 16'hFFFF,
16'h1BB6, 16'hFFFF,
16'h1BB7, 16'hFFFF,
16'h1BB8, 16'hFFFF,
16'h1BB9, 16'hFFFF,
16'h1BBA, 16'hFFFF,
16'h1BBB, 16'hFFFF,
16'h1BBC, 16'hFFFF,
16'h1BBD, 16'hFFFF,
16'h1BBE, 16'hFFFF,
16'h1BBF, 16'hFFFF,
16'h1BC0, 16'hFFFF,
16'h1BC1, 16'hFFFF,
16'h1BC2, 16'hFFFF,
16'h1BC3, 16'hFFFF,
16'h1BC4, 16'hFFFF,
16'h1BC5, 16'hFFFF,
16'h1BC6, 16'hFFFF,
16'h1BC7, 16'hFFFF,
16'h1BC8, 16'hFFFF,
16'h1BC9, 16'hFFFF,
16'h1BCA, 16'hFFFF,
16'h1BCB, 16'hFFFF,
16'h1BCC, 16'hFFFF,
16'h1BCD, 16'hFFFF,
16'h1BCE, 16'hFFFF,
16'h1BCF, 16'hFFFF,
16'h1BD0, 16'hFFFF,
16'h1BD1, 16'hFFFF,
16'h1BD2, 16'hFFFF,
16'h1BD3, 16'hFFFF,
16'h1BD4, 16'hFFFF,
16'h1BD5, 16'hFFFF,
16'h1BD6, 16'hFFFF,
16'h1BD7, 16'hFFFF,
16'h1BD8, 16'hFFFF,
16'h1BD9, 16'hFFFF,
16'h1BDA, 16'hFFFF,
16'h1BDB, 16'hFFFF,
16'h1BDC, 16'hFFFF,
16'h1BDD, 16'hFFFF,
16'h1BDE, 16'hFFFF,
16'h1BDF, 16'hFFFF,
16'h1BE0, 16'hFFFF,
16'h1BE1, 16'hFFFF,
16'h1BE2, 16'hFFFF,
16'h1BE3, 16'hFFFF,
16'h1BE4, 16'hFFFF,
16'h1BE5, 16'hFFFF,
16'h1BE6, 16'hFFFF,
16'h1BE7, 16'hFFFF,
16'h1BE8, 16'hFFFF,
16'h1BE9, 16'hFFFF,
16'h1BEA, 16'hFFFF,
16'h1BEB, 16'hFFFF,
16'h1BEC, 16'hFFFF,
16'h1BED, 16'hFFFF,
16'h1BEE, 16'hFFFF,
16'h1BEF, 16'hFFFF,
16'h1BF0, 16'hFFFF,
16'h1BF1, 16'hFFFF,
16'h1BF2, 16'hFFFF,
16'h1BF3, 16'hFFFF,
16'h1BF4, 16'hFFFF,
16'h1BF5, 16'hFFFF,
16'h1BF6, 16'hFFFF,
16'h1BF7, 16'hFFFF,
16'h1BF8, 16'hFFFF,
16'h1BF9, 16'hFFFF,
16'h1BFA, 16'hFFFF,
16'h1BFB, 16'hFFFF,
16'h1BFC, 16'hFFFF,
16'h1BFD, 16'hFFFF,
16'h1BFE, 16'hFFFF,
16'h1BFF, 16'hFFFF,
16'h1C00, 16'hFFFF,
16'h1C01, 16'hFFFF,
16'h1C02, 16'hFFFF,
16'h1C03, 16'hFFFF,
16'h1C04, 16'hFFFF,
16'h1C05, 16'hFFFF,
16'h1C06, 16'hFFFF,
16'h1C07, 16'hFFFF,
16'h1C08, 16'hFFFF,
16'h1C09, 16'hFFFF,
16'h1C0A, 16'hFFFF,
16'h1C0B, 16'hFFFF,
16'h1C0C, 16'hFFFF,
16'h1C0D, 16'hFFFF,
16'h1C0E, 16'hFFFF,
16'h1C0F, 16'hFFFF,
16'h1C10, 16'hFFFF,
16'h1C11, 16'hFFFF,
16'h1C12, 16'hFFFF,
16'h1C13, 16'hFFFF,
16'h1C14, 16'hFFFF,
16'h1C15, 16'hFFFF,
16'h1C16, 16'hFFFF,
16'h1C17, 16'hFFFF,
16'h1C18, 16'hFFFF,
16'h1C19, 16'hFFFF,
16'h1C1A, 16'hFFFF,
16'h1C1B, 16'hFFFF,
16'h1C1C, 16'hFFFF,
16'h1C1D, 16'hFFFF,
16'h1C1E, 16'hFFFF,
16'h1C1F, 16'hFFFF,
16'h1C20, 16'hFFFF,
16'h1C21, 16'hFFFF,
16'h1C22, 16'hFFFF,
16'h1C23, 16'hFFFF,
16'h1C24, 16'hFFFF,
16'h1C25, 16'hFFFF,
16'h1C26, 16'hFFFF,
16'h1C27, 16'hFFFF,
16'h1C28, 16'hFFFF,
16'h1C29, 16'hFFFF,
16'h1C2A, 16'hFFFF,
16'h1C2B, 16'hFFFF,
16'h1C2C, 16'hFFFF,
16'h1C2D, 16'hFFFF,
16'h1C2E, 16'hFFFF,
16'h1C2F, 16'hFFFF,
16'h1C30, 16'hFFFF,
16'h1C31, 16'hFFFF,
16'h1C32, 16'hFFFF,
16'h1C33, 16'hFFFF,
16'h1C34, 16'hFFFF,
16'h1C35, 16'hFFFF,
16'h1C36, 16'hFFFF,
16'h1C37, 16'hFFFF,
16'h1C38, 16'hFFFF,
16'h1C39, 16'hFFFF,
16'h1C3A, 16'hFFFF,
16'h1C3B, 16'hFFFF,
16'h1C3C, 16'hFFFF,
16'h1C3D, 16'hFFFF,
16'h1C3E, 16'hFFFF,
16'h1C3F, 16'hFFFF,
16'h1C40, 16'hFFFF,
16'h1C41, 16'hFFFF,
16'h1C42, 16'hFFFF,
16'h1C43, 16'hFFFF,
16'h1C44, 16'hFFFF,
16'h1C45, 16'hFFFF,
16'h1C46, 16'hFFFF,
16'h1C47, 16'hFFFF,
16'h1C48, 16'hFFFF,
16'h1C49, 16'hFFFF,
16'h1C4A, 16'hFFFF,
16'h1C4B, 16'hFFFF,
16'h1C4C, 16'hFFFF,
16'h1C4D, 16'hFFFF,
16'h1C4E, 16'hFFFF,
16'h1C4F, 16'hFFFF,
16'h1C50, 16'hFFFF,
16'h1C51, 16'hFFFF,
16'h1C52, 16'hFFFF,
16'h1C53, 16'hFFFF,
16'h1C54, 16'hFFFF,
16'h1C55, 16'hFFFF,
16'h1C56, 16'hFFFF,
16'h1C57, 16'hFFFF,
16'h1C58, 16'hFFFF,
16'h1C59, 16'hFFFF,
16'h1C5A, 16'hFFFF,
16'h1C5B, 16'hFFFF,
16'h1C5C, 16'hFFFF,
16'h1C5D, 16'hFFFF,
16'h1C5E, 16'hFFFF,
16'h1C5F, 16'hFFFF,
16'h1C60, 16'hFFFF,
16'h1C61, 16'hFFFF,
16'h1C62, 16'hFFFF,
16'h1C63, 16'hFFFF,
16'h1C64, 16'hFFFF,
16'h1C65, 16'hFFFF,
16'h1C66, 16'hFFFF,
16'h1C67, 16'hFFFF,
16'h1C68, 16'hFFFF,
16'h1C69, 16'hFFFF,
16'h1C6A, 16'hFFFF,
16'h1C6B, 16'hFFFF,
16'h1C6C, 16'hFFFF,
16'h1C6D, 16'hFFFF,
16'h1C6E, 16'hFFFF,
16'h1C6F, 16'hFFFF,
16'h1C70, 16'hFFFF,
16'h1C71, 16'hFFFF,
16'h1C72, 16'hFFFF,
16'h1C73, 16'hFFFF,
16'h1C74, 16'hFFFF,
16'h1C75, 16'hFFFF,
16'h1C76, 16'hFFFF,
16'h1C77, 16'hFFFF,
16'h1C78, 16'hFFFF,
16'h1C79, 16'hFFFF,
16'h1C7A, 16'hFFFF,
16'h1C7B, 16'hFFFF,
16'h1C7C, 16'hFFFF,
16'h1C7D, 16'hFFFF,
16'h1C7E, 16'hFFFF,
16'h1C7F, 16'hFFFF,
16'h1C80, 16'hFFFF,
16'h1C81, 16'hFFFF,
16'h1C82, 16'hFFFF,
16'h1C83, 16'hFFFF,
16'h1C84, 16'hFFFF,
16'h1C85, 16'hFFFF,
16'h1C86, 16'hFFFF,
16'h1C87, 16'hFFFF,
16'h1C88, 16'hFFFF,
16'h1C89, 16'hFFFF,
16'h1C8A, 16'hFFFF,
16'h1C8B, 16'hFFFF,
16'h1C8C, 16'hFFFF,
16'h1C8D, 16'hFFFF,
16'h1C8E, 16'hFFFF,
16'h1C8F, 16'hFFFF,
16'h1C90, 16'hFFFF,
16'h1C91, 16'hFFFF,
16'h1C92, 16'hFFFF,
16'h1C93, 16'hFFFF,
16'h1C94, 16'hFFFF,
16'h1C95, 16'hFFFF,
16'h1C96, 16'hFFFF,
16'h1C97, 16'hFFFF,
16'h1C98, 16'hFFFF,
16'h1C99, 16'hFFFF,
16'h1C9A, 16'hFFFF,
16'h1C9B, 16'hFFFF,
16'h1C9C, 16'hFFFF,
16'h1C9D, 16'hFFFF,
16'h1C9E, 16'hFFFF,
16'h1C9F, 16'hFFFF,
16'h1CA0, 16'hFFFF,
16'h1CA1, 16'hFFFF,
16'h1CA2, 16'hFFFF,
16'h1CA3, 16'hFFFF,
16'h1CA4, 16'hFFFF,
16'h1CA5, 16'hFFFF,
16'h1CA6, 16'hFFFF,
16'h1CA7, 16'hFFFF,
16'h1CA8, 16'hFFFF,
16'h1CA9, 16'hFFFF,
16'h1CAA, 16'hFFFF,
16'h1CAB, 16'hFFFF,
16'h1CAC, 16'hFFFF,
16'h1CAD, 16'hFFFF,
16'h1CAE, 16'hFFFF,
16'h1CAF, 16'hFFFF,
16'h1CB0, 16'hFFFF,
16'h1CB1, 16'hFFFF,
16'h1CB2, 16'hFFFF,
16'h1CB3, 16'hFFFF,
16'h1CB4, 16'hFFFF,
16'h1CB5, 16'hFFFF,
16'h1CB6, 16'hFFFF,
16'h1CB7, 16'hFFFF,
16'h1CB8, 16'hFFFF,
16'h1CB9, 16'hFFFF,
16'h1CBA, 16'hFFFF,
16'h1CBB, 16'hFFFF,
16'h1CBC, 16'hFFFF,
16'h1CBD, 16'hFFFF,
16'h1CBE, 16'hFFFF,
16'h1CBF, 16'hFFFF,
16'h1CC0, 16'hFFFF,
16'h1CC1, 16'hFFFF,
16'h1CC2, 16'hFFFF,
16'h1CC3, 16'hFFFF,
16'h1CC4, 16'hFFFF,
16'h1CC5, 16'hFFFF,
16'h1CC6, 16'hFFFF,
16'h1CC7, 16'hFFFF,
16'h1CC8, 16'hFFFF,
16'h1CC9, 16'hFFFF,
16'h1CCA, 16'hFFFF,
16'h1CCB, 16'hFFFF,
16'h1CCC, 16'hFFFF,
16'h1CCD, 16'hFFFF,
16'h1CCE, 16'hFFFF,
16'h1CCF, 16'hFFFF,
16'h1CD0, 16'hFFFF,
16'h1CD1, 16'hFFFF,
16'h1CD2, 16'hFFFF,
16'h1CD3, 16'hFFFF,
16'h1CD4, 16'hFFFF,
16'h1CD5, 16'hFFFF,
16'h1CD6, 16'hFFFF,
16'h1CD7, 16'hFFFF,
16'h1CD8, 16'hFFFF,
16'h1CD9, 16'hFFFF,
16'h1CDA, 16'hFFFF,
16'h1CDB, 16'hFFFF,
16'h1CDC, 16'hFFFF,
16'h1CDD, 16'hFFFF,
16'h1CDE, 16'hFFFF,
16'h1CDF, 16'hFFFF,
16'h1CE0, 16'hFFFF,
16'h1CE1, 16'hFFFF,
16'h1CE2, 16'hFFFF,
16'h1CE3, 16'hFFFF,
16'h1CE4, 16'hFFFF,
16'h1CE5, 16'hFFFF,
16'h1CE6, 16'hFFFF,
16'h1CE7, 16'hFFFF,
16'h1CE8, 16'hFFFF,
16'h1CE9, 16'hFFFF,
16'h1CEA, 16'hFFFF,
16'h1CEB, 16'hFFFF,
16'h1CEC, 16'hFFFF,
16'h1CED, 16'hFFFF,
16'h1CEE, 16'hFFFF,
16'h1CEF, 16'hFFFF,
16'h1CF0, 16'hFFFF,
16'h1CF1, 16'hFFFF,
16'h1CF2, 16'hFFFF,
16'h1CF3, 16'hFFFF,
16'h1CF4, 16'hFFFF,
16'h1CF5, 16'hFFFF,
16'h1CF6, 16'hFFFF,
16'h1CF7, 16'hFFFF,
16'h1CF8, 16'hFFFF,
16'h1CF9, 16'hFFFF,
16'h1CFA, 16'hFFFF,
16'h1CFB, 16'hFFFF,
16'h1CFC, 16'hFFFF,
16'h1CFD, 16'hFFFF,
16'h1CFE, 16'hFFFF,
16'h1CFF, 16'hFFFF,
16'h1D00, 16'hFFFF,
16'h1D01, 16'hFFFF,
16'h1D02, 16'hFFFF,
16'h1D03, 16'hFFFF,
16'h1D04, 16'hFFFF,
16'h1D05, 16'hFFFF,
16'h1D06, 16'hFFFF,
16'h1D07, 16'hFFFF,
16'h1D08, 16'hFFFF,
16'h1D09, 16'hFFFF,
16'h1D0A, 16'hFFFF,
16'h1D0B, 16'hFFFF,
16'h1D0C, 16'hFFFF,
16'h1D0D, 16'hFFFF,
16'h1D0E, 16'hFFFF,
16'h1D0F, 16'hFFFF,
16'h1D10, 16'hFFFF,
16'h1D11, 16'hFFFF,
16'h1D12, 16'hFFFF,
16'h1D13, 16'hFFFF,
16'h1D14, 16'hFFFF,
16'h1D15, 16'hFFFF,
16'h1D16, 16'hFFFF,
16'h1D17, 16'hFFFF,
16'h1D18, 16'hFFFF,
16'h1D19, 16'hFFFF,
16'h1D1A, 16'hFFFF,
16'h1D1B, 16'hFFFF,
16'h1D1C, 16'hFFFF,
16'h1D1D, 16'hFFFF,
16'h1D1E, 16'hFFFF,
16'h1D1F, 16'hFFFF,
16'h1D20, 16'hFFFF,
16'h1D21, 16'hFFFF,
16'h1D22, 16'hFFFF,
16'h1D23, 16'hFFFF,
16'h1D24, 16'hFFFF,
16'h1D25, 16'hFFFF,
16'h1D26, 16'hFFFF,
16'h1D27, 16'hFFFF,
16'h1D28, 16'hFFFF,
16'h1D29, 16'hFFFF,
16'h1D2A, 16'hFFFF,
16'h1D2B, 16'hFFFF,
16'h1D2C, 16'hFFFF,
16'h1D2D, 16'hFFFF,
16'h1D2E, 16'hFFFF,
16'h1D2F, 16'hFFFF,
16'h1D30, 16'hFFFF,
16'h1D31, 16'hFFFF,
16'h1D32, 16'hFFFF,
16'h1D33, 16'hFFFF,
16'h1D34, 16'hFFFF,
16'h1D35, 16'hFFFF,
16'h1D36, 16'hFFFF,
16'h1D37, 16'hFFFF,
16'h1D38, 16'hFFFF,
16'h1D39, 16'hFFFF,
16'h1D3A, 16'hFFFF,
16'h1D3B, 16'hFFFF,
16'h1D3C, 16'hFFFF,
16'h1D3D, 16'hFFFF,
16'h1D3E, 16'hFFFF,
16'h1D3F, 16'hFFFF,
16'h1D40, 16'hFFFF,
16'h1D41, 16'hFFFF,
16'h1D42, 16'hFFFF,
16'h1D43, 16'hFFFF,
16'h1D44, 16'hFFFF,
16'h1D45, 16'hFFFF,
16'h1D46, 16'hFFFF,
16'h1D47, 16'hFFFF,
16'h1D48, 16'hFFFF,
16'h1D49, 16'hFFFF,
16'h1D4A, 16'hFFFF,
16'h1D4B, 16'hFFFF,
16'h1D4C, 16'hFFFF,
16'h1D4D, 16'hFFFF,
16'h1D4E, 16'hFFFF,
16'h1D4F, 16'hFFFF,
16'h1D50, 16'hFFFF,
16'h1D51, 16'hFFFF,
16'h1D52, 16'hFFFF,
16'h1D53, 16'hFFFF,
16'h1D54, 16'hFFFF,
16'h1D55, 16'hFFFF,
16'h1D56, 16'hFFFF,
16'h1D57, 16'hFFFF,
16'h1D58, 16'hFFFF,
16'h1D59, 16'hFFFF,
16'h1D5A, 16'hFFFF,
16'h1D5B, 16'hFFFF,
16'h1D5C, 16'hFFFF,
16'h1D5D, 16'hFFFF,
16'h1D5E, 16'hFFFF,
16'h1D5F, 16'hFFFF,
16'h1D60, 16'hFFFF,
16'h1D61, 16'hFFFF,
16'h1D62, 16'hFFFF,
16'h1D63, 16'hFFFF,
16'h1D64, 16'hFFFF,
16'h1D65, 16'hFFFF,
16'h1D66, 16'hFFFF,
16'h1D67, 16'hFFFF,
16'h1D68, 16'hFFFF,
16'h1D69, 16'hFFFF,
16'h1D6A, 16'hFFFF,
16'h1D6B, 16'hFFFF,
16'h1D6C, 16'hFFFF,
16'h1D6D, 16'hFFFF,
16'h1D6E, 16'hFFFF,
16'h1D6F, 16'hFFFF,
16'h1D70, 16'hFFFF,
16'h1D71, 16'hFFFF,
16'h1D72, 16'hFFFF,
16'h1D73, 16'hFFFF,
16'h1D74, 16'hFFFF,
16'h1D75, 16'hFFFF,
16'h1D76, 16'hFFFF,
16'h1D77, 16'hFFFF,
16'h1D78, 16'hFFFF,
16'h1D79, 16'hFFFF,
16'h1D7A, 16'hFFFF,
16'h1D7B, 16'hFFFF,
16'h1D7C, 16'hFFFF,
16'h1D7D, 16'hFFFF,
16'h1D7E, 16'hFFFF,
16'h1D7F, 16'hFFFF,
16'h1D80, 16'hFFFF,
16'h1D81, 16'hFFFF,
16'h1D82, 16'hFFFF,
16'h1D83, 16'hFFFF,
16'h1D84, 16'hFFFF,
16'h1D85, 16'hFFFF,
16'h1D86, 16'hFFFF,
16'h1D87, 16'hFFFF,
16'h1D88, 16'hFFFF,
16'h1D89, 16'hFFFF,
16'h1D8A, 16'hFFFF,
16'h1D8B, 16'hFFFF,
16'h1D8C, 16'hFFFF,
16'h1D8D, 16'hFFFF,
16'h1D8E, 16'hFFFF,
16'h1D8F, 16'hFFFF,
16'h1D90, 16'hFFFF,
16'h1D91, 16'hFFFF,
16'h1D92, 16'hFFFF,
16'h1D93, 16'hFFFF,
16'h1D94, 16'hFFFF,
16'h1D95, 16'hFFFF,
16'h1D96, 16'hFFFF,
16'h1D97, 16'hFFFF,
16'h1D98, 16'hFFFF,
16'h1D99, 16'hFFFF,
16'h1D9A, 16'hFFFF,
16'h1D9B, 16'hFFFF,
16'h1D9C, 16'hFFFF,
16'h1D9D, 16'hFFFF,
16'h1D9E, 16'hFFFF,
16'h1D9F, 16'hFFFF,
16'h1DA0, 16'hFFFF,
16'h1DA1, 16'hFFFF,
16'h1DA2, 16'hFFFF,
16'h1DA3, 16'hFFFF,
16'h1DA4, 16'hFFFF,
16'h1DA5, 16'hFFFF,
16'h1DA6, 16'hFFFF,
16'h1DA7, 16'hFFFF,
16'h1DA8, 16'hFFFF,
16'h1DA9, 16'hFFFF,
16'h1DAA, 16'hFFFF,
16'h1DAB, 16'hFFFF,
16'h1DAC, 16'hFFFF,
16'h1DAD, 16'hFFFF,
16'h1DAE, 16'hFFFF,
16'h1DAF, 16'hFFFF,
16'h1DB0, 16'hFFFF,
16'h1DB1, 16'hFFFF,
16'h1DB2, 16'hFFFF,
16'h1DB3, 16'hFFFF,
16'h1DB4, 16'hFFFF,
16'h1DB5, 16'hFFFF,
16'h1DB6, 16'hFFFF,
16'h1DB7, 16'hFFFF,
16'h1DB8, 16'hFFFF,
16'h1DB9, 16'hFFFF,
16'h1DBA, 16'hFFFF,
16'h1DBB, 16'hFFFF,
16'h1DBC, 16'hFFFF,
16'h1DBD, 16'hFFFF,
16'h1DBE, 16'hFFFF,
16'h1DBF, 16'hFFFF,
16'h1DC0, 16'hFFFF,
16'h1DC1, 16'hFFFF,
16'h1DC2, 16'hFFFF,
16'h1DC3, 16'hFFFF,
16'h1DC4, 16'hFFFF,
16'h1DC5, 16'hFFFF,
16'h1DC6, 16'hFFFF,
16'h1DC7, 16'hFFFF,
16'h1DC8, 16'hFFFF,
16'h1DC9, 16'hFFFF,
16'h1DCA, 16'hFFFF,
16'h1DCB, 16'hFFFF,
16'h1DCC, 16'hFFFF,
16'h1DCD, 16'hFFFF,
16'h1DCE, 16'hFFFF,
16'h1DCF, 16'hFFFF,
16'h1DD0, 16'hFFFF,
16'h1DD1, 16'hFFFF,
16'h1DD2, 16'hFFFF,
16'h1DD3, 16'hFFFF,
16'h1DD4, 16'hFFFF,
16'h1DD5, 16'hFFFF,
16'h1DD6, 16'hFFFF,
16'h1DD7, 16'hFFFF,
16'h1DD8, 16'hFFFF,
16'h1DD9, 16'hFFFF,
16'h1DDA, 16'hFFFF,
16'h1DDB, 16'hFFFF,
16'h1DDC, 16'hFFFF,
16'h1DDD, 16'hFFFF,
16'h1DDE, 16'hFFFF,
16'h1DDF, 16'hFFFF,
16'h1DE0, 16'hFFFF,
16'h1DE1, 16'hFFFF,
16'h1DE2, 16'hFFFF,
16'h1DE3, 16'hFFFF,
16'h1DE4, 16'hFFFF,
16'h1DE5, 16'hFFFF,
16'h1DE6, 16'hFFFF,
16'h1DE7, 16'hFFFF,
16'h1DE8, 16'hFFFF,
16'h1DE9, 16'hFFFF,
16'h1DEA, 16'hFFFF,
16'h1DEB, 16'hFFFF,
16'h1DEC, 16'hFFFF,
16'h1DED, 16'hFFFF,
16'h1DEE, 16'hFFFF,
16'h1DEF, 16'hFFFF,
16'h1DF0, 16'hFFFF,
16'h1DF1, 16'hFFFF,
16'h1DF2, 16'hFFFF,
16'h1DF3, 16'hFFFF,
16'h1DF4, 16'hFFFF,
16'h1DF5, 16'hFFFF,
16'h1DF6, 16'hFFFF,
16'h1DF7, 16'hFFFF,
16'h1DF8, 16'hFFFF,
16'h1DF9, 16'hFFFF,
16'h1DFA, 16'hFFFF,
16'h1DFB, 16'hFFFF,
16'h1DFC, 16'hFFFF,
16'h1DFD, 16'hFFFF,
16'h1DFE, 16'hFFFF,
16'h1DFF, 16'hFFFF,
16'h1E00, 16'hFFFF,
16'h1E01, 16'hFFFF,
16'h1E02, 16'hFFFF,
16'h1E03, 16'hFFFF,
16'h1E04, 16'hFFFF,
16'h1E05, 16'hFFFF,
16'h1E06, 16'hFFFF,
16'h1E07, 16'hFFFF,
16'h1E08, 16'hFFFF,
16'h1E09, 16'hFFFF,
16'h1E0A, 16'hFFFF,
16'h1E0B, 16'hFFFF,
16'h1E0C, 16'hFFFF,
16'h1E0D, 16'hFFFF,
16'h1E0E, 16'hFFFF,
16'h1E0F, 16'hFFFF,
16'h1E10, 16'hFFFF,
16'h1E11, 16'hFFFF,
16'h1E12, 16'hFFFF,
16'h1E13, 16'hFFFF,
16'h1E14, 16'hFFFF,
16'h1E15, 16'hFFFF,
16'h1E16, 16'hFFFF,
16'h1E17, 16'hFFFF,
16'h1E18, 16'hFFFF,
16'h1E19, 16'hFFFF,
16'h1E1A, 16'hFFFF,
16'h1E1B, 16'hFFFF,
16'h1E1C, 16'hFFFF,
16'h1E1D, 16'hFFFF,
16'h1E1E, 16'hFFFF,
16'h1E1F, 16'hFFFF,
16'h1E20, 16'hFFFF,
16'h1E21, 16'hFFFF,
16'h1E22, 16'hFFFF,
16'h1E23, 16'hFFFF,
16'h1E24, 16'hFFFF,
16'h1E25, 16'hFFFF,
16'h1E26, 16'hFFFF,
16'h1E27, 16'hFFFF,
16'h1E28, 16'hFFFF,
16'h1E29, 16'hFFFF,
16'h1E2A, 16'hFFFF,
16'h1E2B, 16'hFFFF,
16'h1E2C, 16'hFFFF,
16'h1E2D, 16'hFFFF,
16'h1E2E, 16'hFFFF,
16'h1E2F, 16'hFFFF,
16'h1E30, 16'hFFFF,
16'h1E31, 16'hFFFF,
16'h1E32, 16'hFFFF,
16'h1E33, 16'hFFFF,
16'h1E34, 16'hFFFF,
16'h1E35, 16'hFFFF,
16'h1E36, 16'hFFFF,
16'h1E37, 16'hFFFF,
16'h1E38, 16'hFFFF,
16'h1E39, 16'hFFFF,
16'h1E3A, 16'hFFFF,
16'h1E3B, 16'hFFFF,
16'h1E3C, 16'hFFFF,
16'h1E3D, 16'hFFFF,
16'h1E3E, 16'hFFFF,
16'h1E3F, 16'hFFFF,
16'h1E40, 16'hFFFF,
16'h1E41, 16'hFFFF,
16'h1E42, 16'hFFFF,
16'h1E43, 16'hFFFF,
16'h1E44, 16'hFFFF,
16'h1E45, 16'hFFFF,
16'h1E46, 16'hFFFF,
16'h1E47, 16'hFFFF,
16'h1E48, 16'hFFFF,
16'h1E49, 16'hFFFF,
16'h1E4A, 16'hFFFF,
16'h1E4B, 16'hFFFF,
16'h1E4C, 16'hFFFF,
16'h1E4D, 16'hFFFF,
16'h1E4E, 16'hFFFF,
16'h1E4F, 16'hFFFF,
16'h1E50, 16'hFFFF,
16'h1E51, 16'hFFFF,
16'h1E52, 16'hFFFF,
16'h1E53, 16'hFFFF,
16'h1E54, 16'hFFFF,
16'h1E55, 16'hFFFF,
16'h1E56, 16'hFFFF,
16'h1E57, 16'hFFFF,
16'h1E58, 16'hFFFF,
16'h1E59, 16'hFFFF,
16'h1E5A, 16'hFFFF,
16'h1E5B, 16'hFFFF,
16'h1E5C, 16'hFFFF,
16'h1E5D, 16'hFFFF,
16'h1E5E, 16'hFFFF,
16'h1E5F, 16'hFFFF,
16'h1E60, 16'hFFFF,
16'h1E61, 16'hFFFF,
16'h1E62, 16'hFFFF,
16'h1E63, 16'hFFFF,
16'h1E64, 16'hFFFF,
16'h1E65, 16'hFFFF,
16'h1E66, 16'hFFFF,
16'h1E67, 16'hFFFF,
16'h1E68, 16'hFFFF,
16'h1E69, 16'hFFFF,
16'h1E6A, 16'hFFFF,
16'h1E6B, 16'hFFFF,
16'h1E6C, 16'hFFFF,
16'h1E6D, 16'hFFFF,
16'h1E6E, 16'hFFFF,
16'h1E6F, 16'hFFFF,
16'h1E70, 16'hFFFF,
16'h1E71, 16'hFFFF,
16'h1E72, 16'hFFFF,
16'h1E73, 16'hFFFF,
16'h1E74, 16'hFFFF,
16'h1E75, 16'hFFFF,
16'h1E76, 16'hFFFF,
16'h1E77, 16'hFFFF,
16'h1E78, 16'hFFFF,
16'h1E79, 16'hFFFF,
16'h1E7A, 16'hFFFF,
16'h1E7B, 16'hFFFF,
16'h1E7C, 16'hFFFF,
16'h1E7D, 16'hFFFF,
16'h1E7E, 16'hFFFF,
16'h1E7F, 16'hFFFF,
16'h1E80, 16'hFFFF,
16'h1E81, 16'hFFFF,
16'h1E82, 16'hFFFF,
16'h1E83, 16'hFFFF,
16'h1E84, 16'hFFFF,
16'h1E85, 16'hFFFF,
16'h1E86, 16'hFFFF,
16'h1E87, 16'hFFFF,
16'h1E88, 16'hFFFF,
16'h1E89, 16'hFFFF,
16'h1E8A, 16'hFFFF,
16'h1E8B, 16'hFFFF,
16'h1E8C, 16'hFFFF,
16'h1E8D, 16'hFFFF,
16'h1E8E, 16'hFFFF,
16'h1E8F, 16'hFFFF,
16'h1E90, 16'hFFFF,
16'h1E91, 16'hFFFF,
16'h1E92, 16'hFFFF,
16'h1E93, 16'hFFFF,
16'h1E94, 16'hFFFF,
16'h1E95, 16'hFFFF,
16'h1E96, 16'hFFFF,
16'h1E97, 16'hFFFF,
16'h1E98, 16'hFFFF,
16'h1E99, 16'hFFFF,
16'h1E9A, 16'hFFFF,
16'h1E9B, 16'hFFFF,
16'h1E9C, 16'hFFFF,
16'h1E9D, 16'hFFFF,
16'h1E9E, 16'hFFFF,
16'h1E9F, 16'hFFFF,
16'h1EA0, 16'hFFFF,
16'h1EA1, 16'hFFFF,
16'h1EA2, 16'hFFFF,
16'h1EA3, 16'hFFFF,
16'h1EA4, 16'hFFFF,
16'h1EA5, 16'hFFFF,
16'h1EA6, 16'hFFFF,
16'h1EA7, 16'hFFFF,
16'h1EA8, 16'hFFFF,
16'h1EA9, 16'hFFFF,
16'h1EAA, 16'hFFFF,
16'h1EAB, 16'hFFFF,
16'h1EAC, 16'hFFFF,
16'h1EAD, 16'hFFFF,
16'h1EAE, 16'hFFFF,
16'h1EAF, 16'hFFFF,
16'h1EB0, 16'hFFFF,
16'h1EB1, 16'hFFFF,
16'h1EB2, 16'hFFFF,
16'h1EB3, 16'hFFFF,
16'h1EB4, 16'hFFFF,
16'h1EB5, 16'hFFFF,
16'h1EB6, 16'hFFFF,
16'h1EB7, 16'hFFFF,
16'h1EB8, 16'hFFFF,
16'h1EB9, 16'hFFFF,
16'h1EBA, 16'hFFFF,
16'h1EBB, 16'hFFFF,
16'h1EBC, 16'hFFFF,
16'h1EBD, 16'hFFFF,
16'h1EBE, 16'hFFFF,
16'h1EBF, 16'hFFFF,
16'h1EC0, 16'hFFFF,
16'h1EC1, 16'hFFFF,
16'h1EC2, 16'hFFFF,
16'h1EC3, 16'hFFFF,
16'h1EC4, 16'hFFFF,
16'h1EC5, 16'hFFFF,
16'h1EC6, 16'hFFFF,
16'h1EC7, 16'hFFFF,
16'h1EC8, 16'hFFFF,
16'h1EC9, 16'hFFFF,
16'h1ECA, 16'hFFFF,
16'h1ECB, 16'hFFFF,
16'h1ECC, 16'hFFFF,
16'h1ECD, 16'hFFFF,
16'h1ECE, 16'hFFFF,
16'h1ECF, 16'hFFFF,
16'h1ED0, 16'hFFFF,
16'h1ED1, 16'hFFFF,
16'h1ED2, 16'hFFFF,
16'h1ED3, 16'hFFFF,
16'h1ED4, 16'hFFFF,
16'h1ED5, 16'hFFFF,
16'h1ED6, 16'hFFFF,
16'h1ED7, 16'hFFFF,
16'h1ED8, 16'hFFFF,
16'h1ED9, 16'hFFFF,
16'h1EDA, 16'hFFFF,
16'h1EDB, 16'hFFFF,
16'h1EDC, 16'hFFFF,
16'h1EDD, 16'hFFFF,
16'h1EDE, 16'hFFFF,
16'h1EDF, 16'hFFFF,
16'h1EE0, 16'hFFFF,
16'h1EE1, 16'hFFFF,
16'h1EE2, 16'hFFFF,
16'h1EE3, 16'hFFFF,
16'h1EE4, 16'hFFFF,
16'h1EE5, 16'hFFFF,
16'h1EE6, 16'hFFFF,
16'h1EE7, 16'hFFFF,
16'h1EE8, 16'hFFFF,
16'h1EE9, 16'hFFFF,
16'h1EEA, 16'hFFFF,
16'h1EEB, 16'hFFFF,
16'h1EEC, 16'hFFFF,
16'h1EED, 16'hFFFF,
16'h1EEE, 16'hFFFF,
16'h1EEF, 16'hFFFF,
16'h1EF0, 16'hFFFF,
16'h1EF1, 16'hFFFF,
16'h1EF2, 16'hFFFF,
16'h1EF3, 16'hFFFF,
16'h1EF4, 16'hFFFF,
16'h1EF5, 16'hFFFF,
16'h1EF6, 16'hFFFF,
16'h1EF7, 16'hFFFF,
16'h1EF8, 16'hFFFF,
16'h1EF9, 16'hFFFF,
16'h1EFA, 16'hFFFF,
16'h1EFB, 16'hFFFF,
16'h1EFC, 16'hFFFF,
16'h1EFD, 16'hFFFF,
16'h1EFE, 16'hFFFF,
16'h1EFF, 16'hFFFF,
16'h1F00, 16'hFFFF,
16'h1F01, 16'hFFFF,
16'h1F02, 16'hFFFF,
16'h1F03, 16'hFFFF,
16'h1F04, 16'hFFFF,
16'h1F05, 16'hFFFF,
16'h1F06, 16'hFFFF,
16'h1F07, 16'hFFFF,
16'h1F08, 16'hFFFF,
16'h1F09, 16'hFFFF,
16'h1F0A, 16'hFFFF,
16'h1F0B, 16'hFFFF,
16'h1F0C, 16'hFFFF,
16'h1F0D, 16'hFFFF,
16'h1F0E, 16'hFFFF,
16'h1F0F, 16'hFFFF,
16'h1F10, 16'hFFFF,
16'h1F11, 16'hFFFF,
16'h1F12, 16'hFFFF,
16'h1F13, 16'hFFFF,
16'h1F14, 16'hFFFF,
16'h1F15, 16'hFFFF,
16'h1F16, 16'hFFFF,
16'h1F17, 16'hFFFF,
16'h1F18, 16'hFFFF,
16'h1F19, 16'hFFFF,
16'h1F1A, 16'hFFFF,
16'h1F1B, 16'hFFFF,
16'h1F1C, 16'hFFFF,
16'h1F1D, 16'hFFFF,
16'h1F1E, 16'hFFFF,
16'h1F1F, 16'hFFFF,
16'h1F20, 16'hFFFF,
16'h1F21, 16'hFFFF,
16'h1F22, 16'hFFFF,
16'h1F23, 16'hFFFF,
16'h1F24, 16'hFFFF,
16'h1F25, 16'hFFFF,
16'h1F26, 16'hFFFF,
16'h1F27, 16'hFFFF,
16'h1F28, 16'hFFFF,
16'h1F29, 16'hFFFF,
16'h1F2A, 16'hFFFF,
16'h1F2B, 16'hFFFF,
16'h1F2C, 16'hFFFF,
16'h1F2D, 16'hFFFF,
16'h1F2E, 16'hFFFF,
16'h1F2F, 16'hFFFF,
16'h1F30, 16'hFFFF,
16'h1F31, 16'hFFFF,
16'h1F32, 16'hFFFF,
16'h1F33, 16'hFFFF,
16'h1F34, 16'hFFFF,
16'h1F35, 16'hFFFF,
16'h1F36, 16'hFFFF,
16'h1F37, 16'hFFFF,
16'h1F38, 16'hFFFF,
16'h1F39, 16'hFFFF,
16'h1F3A, 16'hFFFF,
16'h1F3B, 16'hFFFF,
16'h1F3C, 16'hFFFF,
16'h1F3D, 16'hFFFF,
16'h1F3E, 16'hFFFF,
16'h1F3F, 16'hFFFF,
16'h1F40, 16'hFFFF,
16'h1F41, 16'hFFFF,
16'h1F42, 16'hFFFF,
16'h1F43, 16'hFFFF,
16'h1F44, 16'hFFFF,
16'h1F45, 16'hFFFF,
16'h1F46, 16'hFFFF,
16'h1F47, 16'hFFFF,
16'h1F48, 16'hFFFF,
16'h1F49, 16'hFFFF,
16'h1F4A, 16'hFFFF,
16'h1F4B, 16'hFFFF,
16'h1F4C, 16'hFFFF,
16'h1F4D, 16'hFFFF,
16'h1F4E, 16'hFFFF,
16'h1F4F, 16'hFFFF,
16'h1F50, 16'hFFFF,
16'h1F51, 16'hFFFF,
16'h1F52, 16'hFFFF,
16'h1F53, 16'hFFFF,
16'h1F54, 16'hFFFF,
16'h1F55, 16'hFFFF,
16'h1F56, 16'hFFFF,
16'h1F57, 16'hFFFF,
16'h1F58, 16'hFFFF,
16'h1F59, 16'hFFFF,
16'h1F5A, 16'hFFFF,
16'h1F5B, 16'hFFFF,
16'h1F5C, 16'hFFFF,
16'h1F5D, 16'hFFFF,
16'h1F5E, 16'hFFFF,
16'h1F5F, 16'hFFFF,
16'h1F60, 16'hFFFF,
16'h1F61, 16'hFFFF,
16'h1F62, 16'hFFFF,
16'h1F63, 16'hFFFF,
16'h1F64, 16'hFFFF,
16'h1F65, 16'hFFFF,
16'h1F66, 16'hFFFF,
16'h1F67, 16'hFFFF,
16'h1F68, 16'hFFFF,
16'h1F69, 16'hFFFF,
16'h1F6A, 16'hFFFF,
16'h1F6B, 16'hFFFF,
16'h1F6C, 16'hFFFF,
16'h1F6D, 16'hFFFF,
16'h1F6E, 16'hFFFF,
16'h1F6F, 16'hFFFF,
16'h1F70, 16'hFFFF,
16'h1F71, 16'hFFFF,
16'h1F72, 16'hFFFF,
16'h1F73, 16'hFFFF,
16'h1F74, 16'hFFFF,
16'h1F75, 16'hFFFF,
16'h1F76, 16'hFFFF,
16'h1F77, 16'hFFFF,
16'h1F78, 16'hFFFF,
16'h1F79, 16'hFFFF,
16'h1F7A, 16'hFFFF,
16'h1F7B, 16'hFFFF,
16'h1F7C, 16'hFFFF,
16'h1F7D, 16'hFFFF,
16'h1F7E, 16'hFFFF,
16'h1F7F, 16'hFFFF,
16'h1F80, 16'hFFFF,
16'h1F81, 16'hFFFF,
16'h1F82, 16'hFFFF,
16'h1F83, 16'hFFFF,
16'h1F84, 16'hFFFF,
16'h1F85, 16'hFFFF,
16'h1F86, 16'hFFFF,
16'h1F87, 16'hFFFF,
16'h1F88, 16'hFFFF,
16'h1F89, 16'hFFFF,
16'h1F8A, 16'hFFFF,
16'h1F8B, 16'hFFFF,
16'h1F8C, 16'hFFFF,
16'h1F8D, 16'hFFFF,
16'h1F8E, 16'hFFFF,
16'h1F8F, 16'hFFFF,
16'h1F90, 16'hFFFF,
16'h1F91, 16'hFFFF,
16'h1F92, 16'hFFFF,
16'h1F93, 16'hFFFF,
16'h1F94, 16'hFFFF,
16'h1F95, 16'hFFFF,
16'h1F96, 16'hFFFF,
16'h1F97, 16'hFFFF,
16'h1F98, 16'hFFFF,
16'h1F99, 16'hFFFF,
16'h1F9A, 16'hFFFF,
16'h1F9B, 16'hFFFF,
16'h1F9C, 16'hFFFF,
16'h1F9D, 16'hFFFF,
16'h1F9E, 16'hFFFF,
16'h1F9F, 16'hFFFF,
16'h1FA0, 16'hFFFF,
16'h1FA1, 16'hFFFF,
16'h1FA2, 16'hFFFF,
16'h1FA3, 16'hFFFF,
16'h1FA4, 16'hFFFF,
16'h1FA5, 16'hFFFF,
16'h1FA6, 16'hFFFF,
16'h1FA7, 16'hFFFF,
16'h1FA8, 16'hFFFF,
16'h1FA9, 16'hFFFF,
16'h1FAA, 16'hFFFF,
16'h1FAB, 16'hFFFF,
16'h1FAC, 16'hFFFF,
16'h1FAD, 16'hFFFF,
16'h1FAE, 16'hFFFF,
16'h1FAF, 16'hFFFF,
16'h1FB0, 16'hFFFF,
16'h1FB1, 16'hFFFF,
16'h1FB2, 16'hFFFF,
16'h1FB3, 16'hFFFF,
16'h1FB4, 16'hFFFF,
16'h1FB5, 16'hFFFF,
16'h1FB6, 16'hFFFF,
16'h1FB7, 16'hFFFF,
16'h1FB8, 16'hFFFF,
16'h1FB9, 16'hFFFF,
16'h1FBA, 16'hFFFF,
16'h1FBB, 16'hFFFF,
16'h1FBC, 16'hFFFF,
16'h1FBD, 16'hFFFF,
16'h1FBE, 16'hFFFF,
16'h1FBF, 16'hFFFF,
16'h1FC0, 16'hFFFF,
16'h1FC1, 16'hFFFF,
16'h1FC2, 16'hFFFF,
16'h1FC3, 16'hFFFF,
16'h1FC4, 16'hFFFF,
16'h1FC5, 16'hFFFF,
16'h1FC6, 16'hFFFF,
16'h1FC7, 16'hFFFF,
16'h1FC8, 16'hFFFF,
16'h1FC9, 16'hFFFF,
16'h1FCA, 16'hFFFF,
16'h1FCB, 16'hFFFF,
16'h1FCC, 16'hFFFF,
16'h1FCD, 16'hFFFF,
16'h1FCE, 16'hFFFF,
16'h1FCF, 16'hFFFF,
16'h1FD0, 16'hFFFF,
16'h1FD1, 16'hFFFF,
16'h1FD2, 16'hFFFF,
16'h1FD3, 16'hFFFF,
16'h1FD4, 16'hFFFF,
16'h1FD5, 16'hFFFF,
16'h1FD6, 16'hFFFF,
16'h1FD7, 16'hFFFF,
16'h1FD8, 16'hFFFF,
16'h1FD9, 16'hFFFF,
16'h1FDA, 16'hFFFF,
16'h1FDB, 16'hFFFF,
16'h1FDC, 16'hFFFF,
16'h1FDD, 16'hFFFF,
16'h1FDE, 16'hFFFF,
16'h1FDF, 16'hFFFF,
16'h1FE0, 16'hFFFF,
16'h1FE1, 16'hFFFF,
16'h1FE2, 16'hFFFF,
16'h1FE3, 16'hFFFF,
16'h1FE4, 16'hFFFF,
16'h1FE5, 16'hFFFF,
16'h1FE6, 16'hFFFF,
16'h1FE7, 16'hFFFF,
16'h1FE8, 16'hFFFF,
16'h1FE9, 16'hFFFF,
16'h1FEA, 16'hFFFF,
16'h1FEB, 16'hFFFF,
16'h1FEC, 16'hFFFF,
16'h1FED, 16'hFFFF,
16'h1FEE, 16'hFFFF,
16'h1FEF, 16'hFFFF,
16'h1FF0, 16'hFFFF,
16'h1FF1, 16'hFFFF,
16'h1FF2, 16'hFFFF,
16'h1FF3, 16'hFFFF,
16'h1FF4, 16'hFFFF,
16'h1FF5, 16'hFFFF,
16'h1FF6, 16'hFFFF,
16'h1FF7, 16'hFFFF,
16'h1FF8, 16'hFFFF,
16'h1FF9, 16'hFFFF,
16'h1FFA, 16'hFFFF,
16'h1FFB, 16'hFFFF,
16'h1FFC, 16'hFFFF,
16'h1FFD, 16'hFFFF,
16'h1FFE, 16'hFFFF,
16'h1FFF, 16'hFFFF,
16'h2000, 16'h0000,
16'h2001, 16'h0000,
16'h2002, 16'h0000,
16'h2003, 16'h0000,
16'h2004, 16'h0000,
16'h2005, 16'h0000,
16'h2006, 16'h0000,
16'h2007, 16'h0000,
16'h2008, 16'h0000,
16'h2009, 16'h0000,
16'h200A, 16'h0000,
16'h200B, 16'h0000,
16'h200C, 16'h0000,
16'h200D, 16'h0000,
16'h200E, 16'h0000,
16'h200F, 16'h0000,
16'h2010, 16'h0000,
16'h2011, 16'h0000,
16'h2012, 16'h0000,
16'h2013, 16'h0000,
16'h2014, 16'h0000,
16'h2015, 16'h0000,
16'h2016, 16'h0000,
16'h2017, 16'h0000,
16'h2018, 16'h0000,
16'h2019, 16'h0000,
16'h201A, 16'h0000,
16'h201B, 16'h0000,
16'h201C, 16'h0000,
16'h201D, 16'h0000,
16'h201E, 16'h0000,
16'h201F, 16'h0000,
16'h2020, 16'h0000,
16'h2021, 16'h0000,
16'h2022, 16'h0000,
16'h2023, 16'h0000,
16'h2024, 16'h0000,
16'h2025, 16'h0000,
16'h2026, 16'h0000,
16'h2027, 16'h0000,
16'h2028, 16'h0000,
16'h2029, 16'h0000,
16'h202A, 16'h0000,
16'h202B, 16'h0000,
16'h202C, 16'h0000,
16'h202D, 16'h0000,
16'h202E, 16'h0000,
16'h202F, 16'h0000,
16'h2030, 16'h0000,
16'h2031, 16'h0000,
16'h2032, 16'h0000,
16'h2033, 16'h0000,
16'h2034, 16'h0000,
16'h2035, 16'h0000,
16'h2036, 16'h0000,
16'h2037, 16'h0000,
16'h2038, 16'h0000,
16'h2039, 16'h0000,
16'h203A, 16'h0000,
16'h203B, 16'h0000,
16'h203C, 16'h0000,
16'h203D, 16'h0000,
16'h203E, 16'h0000,
16'h203F, 16'h0000,
16'h2040, 16'h0000,
16'h2041, 16'h0000,
16'h2042, 16'h0000,
16'h2043, 16'h0000,
16'h2044, 16'h0000,
16'h2045, 16'h0000,
16'h2046, 16'h0000,
16'h2047, 16'h0000,
16'h2048, 16'h0000,
16'h2049, 16'h0000,
16'h204A, 16'h0000,
16'h204B, 16'h0000,
16'h204C, 16'h0000,
16'h204D, 16'h0000,
16'h204E, 16'h0000,
16'h204F, 16'h0000,
16'h2050, 16'h0000,
16'h2051, 16'h0000,
16'h2052, 16'h0000,
16'h2053, 16'h0000,
16'h2054, 16'h0000,
16'h2055, 16'h0000,
16'h2056, 16'h0000,
16'h2057, 16'h0000,
16'h2058, 16'h0000,
16'h2059, 16'h0000,
16'h205A, 16'h0000,
16'h205B, 16'h0000,
16'h205C, 16'h0000,
16'h205D, 16'h0000,
16'h205E, 16'h0000,
16'h205F, 16'h0000,
16'h2060, 16'h0000,
16'h2061, 16'h0000,
16'h2062, 16'h0000,
16'h2063, 16'h0000,
16'h2064, 16'h0000,
16'h2065, 16'h0000,
16'h2066, 16'h0000,
16'h2067, 16'h0000,
16'h2068, 16'h0000,
16'h2069, 16'h0000,
16'h206A, 16'h0000,
16'h206B, 16'h0000,
16'h206C, 16'h0000,
16'h206D, 16'h0000,
16'h206E, 16'h0000,
16'h206F, 16'h0000,
16'h2070, 16'h0000,
16'h2071, 16'h0000,
16'h2072, 16'h0000,
16'h2073, 16'h0000,
16'h2074, 16'h0000,
16'h2075, 16'h0000,
16'h2076, 16'h0000,
16'h2077, 16'h0000,
16'h2078, 16'h0000,
16'h2079, 16'h0000,
16'h207A, 16'h0000,
16'h207B, 16'h0000,
16'h207C, 16'h0000,
16'h207D, 16'h0000,
16'h207E, 16'h0000,
16'h207F, 16'h0000,
16'h2080, 16'h0000,
16'h2081, 16'h0000,
16'h2082, 16'h0000,
16'h2083, 16'h0000,
16'h2084, 16'h0000,
16'h2085, 16'h0000,
16'h2086, 16'h0000,
16'h2087, 16'h0000,
16'h2088, 16'h0000,
16'h2089, 16'h0000,
16'h208A, 16'h0000,
16'h208B, 16'h0000,
16'h208C, 16'h0000,
16'h208D, 16'h0000,
16'h208E, 16'h0000,
16'h208F, 16'h0000,
16'h2090, 16'h0000,
16'h2091, 16'h0000,
16'h2092, 16'h0000,
16'h2093, 16'h0000,
16'h2094, 16'h0000,
16'h2095, 16'h0000,
16'h2096, 16'h0000,
16'h2097, 16'h0000,
16'h2098, 16'h0000,
16'h2099, 16'h0000,
16'h209A, 16'h0000,
16'h209B, 16'h0000,
16'h209C, 16'h0000,
16'h209D, 16'h0000,
16'h209E, 16'h0000,
16'h209F, 16'h0000,
16'h20A0, 16'h0000,
16'h20A1, 16'h0000,
16'h20A2, 16'h0000,
16'h20A3, 16'h0000,
16'h20A4, 16'h0000,
16'h20A5, 16'h0000,
16'h20A6, 16'h0000,
16'h20A7, 16'h0000,
16'h20A8, 16'h0000,
16'h20A9, 16'h0000,
16'h20AA, 16'h0000,
16'h20AB, 16'h0000,
16'h20AC, 16'h0000,
16'h20AD, 16'h0000,
16'h20AE, 16'h0000,
16'h20AF, 16'h0000,
16'h20B0, 16'h0000,
16'h20B1, 16'h0000,
16'h20B2, 16'h0000,
16'h20B3, 16'h0000,
16'h20B4, 16'h0000,
16'h20B5, 16'h0000,
16'h20B6, 16'h0000,
16'h20B7, 16'h0000,
16'h20B8, 16'h0000,
16'h20B9, 16'h0000,
16'h20BA, 16'h0000,
16'h20BB, 16'h0000,
16'h20BC, 16'h0000,
16'h20BD, 16'h0000,
16'h20BE, 16'h0000,
16'h20BF, 16'h0000,
16'h20C0, 16'h0000,
16'h20C1, 16'h0000,
16'h20C2, 16'h0000,
16'h20C3, 16'h0000,
16'h20C4, 16'h0000,
16'h20C5, 16'h0000,
16'h20C6, 16'h0000,
16'h20C7, 16'h0000,
16'h20C8, 16'h0000,
16'h20C9, 16'h0000,
16'h20CA, 16'h0000,
16'h20CB, 16'h0000,
16'h20CC, 16'h0000,
16'h20CD, 16'h0000,
16'h20CE, 16'h0000,
16'h20CF, 16'h0000,
16'h20D0, 16'h0000,
16'h20D1, 16'h0000,
16'h20D2, 16'h0000,
16'h20D3, 16'h0000,
16'h20D4, 16'h0000,
16'h20D5, 16'h0000,
16'h20D6, 16'h0000,
16'h20D7, 16'h0000,
16'h20D8, 16'h0000,
16'h20D9, 16'h0000,
16'h20DA, 16'h0000,
16'h20DB, 16'h0000,
16'h20DC, 16'h0000,
16'h20DD, 16'h0000,
16'h20DE, 16'h0000,
16'h20DF, 16'h0000,
16'h20E0, 16'h0000,
16'h20E1, 16'h0000,
16'h20E2, 16'h0000,
16'h20E3, 16'h0000,
16'h20E4, 16'h0000,
16'h20E5, 16'h0000,
16'h20E6, 16'h0000,
16'h20E7, 16'h0000,
16'h20E8, 16'h0000,
16'h20E9, 16'h0000,
16'h20EA, 16'h0000,
16'h20EB, 16'h0000,
16'h20EC, 16'h0000,
16'h20ED, 16'h0000,
16'h20EE, 16'h0000,
16'h20EF, 16'h0000,
16'h20F0, 16'h0000,
16'h20F1, 16'h0000,
16'h20F2, 16'h0000,
16'h20F3, 16'h0000,
16'h20F4, 16'h0000,
16'h20F5, 16'h0000,
16'h20F6, 16'h0000,
16'h20F7, 16'h0000,
16'h20F8, 16'h0000,
16'h20F9, 16'h0000,
16'h20FA, 16'h0000,
16'h20FB, 16'h0000,
16'h20FC, 16'h0000,
16'h20FD, 16'h0000,
16'h20FE, 16'h0000,
16'h20FF, 16'h0000,
16'h2100, 16'h0000,
16'h2101, 16'h0000,
16'h2102, 16'h0000,
16'h2103, 16'h0000,
16'h2104, 16'h0000,
16'h2105, 16'h0000,
16'h2106, 16'h0000,
16'h2107, 16'h0000,
16'h2108, 16'h0000,
16'h2109, 16'h0000,
16'h210A, 16'h0000,
16'h210B, 16'h0000,
16'h210C, 16'h0000,
16'h210D, 16'h0000,
16'h210E, 16'h0000,
16'h210F, 16'h0000,
16'h2110, 16'h0000,
16'h2111, 16'h0000,
16'h2112, 16'h0000,
16'h2113, 16'h0000,
16'h2114, 16'h0000,
16'h2115, 16'h0000,
16'h2116, 16'h0000,
16'h2117, 16'h0000,
16'h2118, 16'h0000,
16'h2119, 16'h0000,
16'h211A, 16'h0000,
16'h211B, 16'h0000,
16'h211C, 16'h0000,
16'h211D, 16'h0000,
16'h211E, 16'h0000,
16'h211F, 16'h0000,
16'h2120, 16'h0000,
16'h2121, 16'h0000,
16'h2122, 16'h0000,
16'h2123, 16'h0000,
16'h2124, 16'h0000,
16'h2125, 16'h0000,
16'h2126, 16'h0000,
16'h2127, 16'h0000,
16'h2128, 16'h0000,
16'h2129, 16'h0000,
16'h212A, 16'h0000,
16'h212B, 16'h0000,
16'h212C, 16'h0000,
16'h212D, 16'h0000,
16'h212E, 16'h0000,
16'h212F, 16'h0000,
16'h2130, 16'h0000,
16'h2131, 16'h0000,
16'h2132, 16'h0000,
16'h2133, 16'h0000,
16'h2134, 16'h0000,
16'h2135, 16'h0000,
16'h2136, 16'h0000,
16'h2137, 16'h0000,
16'h2138, 16'h0000,
16'h2139, 16'h0000,
16'h213A, 16'h0000,
16'h213B, 16'h0000,
16'h213C, 16'h0000,
16'h213D, 16'h0000,
16'h213E, 16'h0000,
16'h213F, 16'h0000,
16'h2140, 16'h0000,
16'h2141, 16'h0000,
16'h2142, 16'h0000,
16'h2143, 16'h0000,
16'h2144, 16'h0000,
16'h2145, 16'h0000,
16'h2146, 16'h0000,
16'h2147, 16'h0000,
16'h2148, 16'h0000,
16'h2149, 16'h0000,
16'h214A, 16'h0000,
16'h214B, 16'h0000,
16'h214C, 16'h0000,
16'h214D, 16'h0000,
16'h214E, 16'h0000,
16'h214F, 16'h0000,
16'h2150, 16'h0000,
16'h2151, 16'h0000,
16'h2152, 16'h0000,
16'h2153, 16'h0000,
16'h2154, 16'h0000,
16'h2155, 16'h0000,
16'h2156, 16'h0000,
16'h2157, 16'h0000,
16'h2158, 16'h0000,
16'h2159, 16'h0000,
16'h215A, 16'h0000,
16'h215B, 16'h0000,
16'h215C, 16'h0000,
16'h215D, 16'h0000,
16'h215E, 16'h0000,
16'h215F, 16'h0000,
16'h2160, 16'h0000,
16'h2161, 16'h0000,
16'h2162, 16'h0000,
16'h2163, 16'h0000,
16'h2164, 16'h0000,
16'h2165, 16'h0000,
16'h2166, 16'h0000,
16'h2167, 16'h0000,
16'h2168, 16'h0000,
16'h2169, 16'h0000,
16'h216A, 16'h0000,
16'h216B, 16'h0000,
16'h216C, 16'h0000,
16'h216D, 16'h0000,
16'h216E, 16'h0000,
16'h216F, 16'h0000,
16'h2170, 16'h0000,
16'h2171, 16'h0000,
16'h2172, 16'h0000,
16'h2173, 16'h0000,
16'h2174, 16'h0000,
16'h2175, 16'h0000,
16'h2176, 16'h0000,
16'h2177, 16'h0000,
16'h2178, 16'h0000,
16'h2179, 16'h0000,
16'h217A, 16'h0000,
16'h217B, 16'h0000,
16'h217C, 16'h0000,
16'h217D, 16'h0000,
16'h217E, 16'h0000,
16'h217F, 16'h0000,
16'h2180, 16'h0000,
16'h2181, 16'h0000,
16'h2182, 16'h0000,
16'h2183, 16'h0000,
16'h2184, 16'h0000,
16'h2185, 16'h0000,
16'h2186, 16'h0000,
16'h2187, 16'h0000,
16'h2188, 16'h0000,
16'h2189, 16'h0000,
16'h218A, 16'h0000,
16'h218B, 16'h0000,
16'h218C, 16'h0000,
16'h218D, 16'h0000,
16'h218E, 16'h0000,
16'h218F, 16'h0000,
16'h2190, 16'h0000,
16'h2191, 16'h0000,
16'h2192, 16'h0000,
16'h2193, 16'h0000,
16'h2194, 16'h0000,
16'h2195, 16'h0000,
16'h2196, 16'h0000,
16'h2197, 16'h0000,
16'h2198, 16'h0000,
16'h2199, 16'h0000,
16'h219A, 16'h0000,
16'h219B, 16'h0000,
16'h219C, 16'h0000,
16'h219D, 16'h0000,
16'h219E, 16'h0000,
16'h219F, 16'h0000,
16'h21A0, 16'h0000,
16'h21A1, 16'h0000,
16'h21A2, 16'h0000,
16'h21A3, 16'h0000,
16'h21A4, 16'h0000,
16'h21A5, 16'h0000,
16'h21A6, 16'h0000,
16'h21A7, 16'h0000,
16'h21A8, 16'h0000,
16'h21A9, 16'h0000,
16'h21AA, 16'h0000,
16'h21AB, 16'h0000,
16'h21AC, 16'h0000,
16'h21AD, 16'h0000,
16'h21AE, 16'h0000,
16'h21AF, 16'h0000,
16'h21B0, 16'h0000,
16'h21B1, 16'h0000,
16'h21B2, 16'h0000,
16'h21B3, 16'h0000,
16'h21B4, 16'h0000,
16'h21B5, 16'h0000,
16'h21B6, 16'h0000,
16'h21B7, 16'h0000,
16'h21B8, 16'h0000,
16'h21B9, 16'h0000,
16'h21BA, 16'h0000,
16'h21BB, 16'h0000,
16'h21BC, 16'h0000,
16'h21BD, 16'h0000,
16'h21BE, 16'h0000,
16'h21BF, 16'h0000,
16'h21C0, 16'h0000,
16'h21C1, 16'h0000,
16'h21C2, 16'h0000,
16'h21C3, 16'h0000,
16'h21C4, 16'h0000,
16'h21C5, 16'h0000,
16'h21C6, 16'h0000,
16'h21C7, 16'h0000,
16'h21C8, 16'h0000,
16'h21C9, 16'h0000,
16'h21CA, 16'h0000,
16'h21CB, 16'h0000,
16'h21CC, 16'h0000,
16'h21CD, 16'h0000,
16'h21CE, 16'h0000,
16'h21CF, 16'h0000,
16'h21D0, 16'h0000,
16'h21D1, 16'h0000,
16'h21D2, 16'h0000,
16'h21D3, 16'h0000,
16'h21D4, 16'h0000,
16'h21D5, 16'h0000,
16'h21D6, 16'h0000,
16'h21D7, 16'h0000,
16'h21D8, 16'h0000,
16'h21D9, 16'h0000,
16'h21DA, 16'h0000,
16'h21DB, 16'h0000,
16'h21DC, 16'h0000,
16'h21DD, 16'h0000,
16'h21DE, 16'h0000,
16'h21DF, 16'h0000,
16'h21E0, 16'h0000,
16'h21E1, 16'h0000,
16'h21E2, 16'h0000,
16'h21E3, 16'h0000,
16'h21E4, 16'h0000,
16'h21E5, 16'h0000,
16'h21E6, 16'h0000,
16'h21E7, 16'h0000,
16'h21E8, 16'h0000,
16'h21E9, 16'h0000,
16'h21EA, 16'h0000,
16'h21EB, 16'h0000,
16'h21EC, 16'h0000,
16'h21ED, 16'h0000,
16'h21EE, 16'h0000,
16'h21EF, 16'h0000,
16'h21F0, 16'h0000,
16'h21F1, 16'h0000,
16'h21F2, 16'h0000,
16'h21F3, 16'h0000,
16'h21F4, 16'h0000,
16'h21F5, 16'h0000,
16'h21F6, 16'h0000,
16'h21F7, 16'h0000,
16'h21F8, 16'h0000,
16'h21F9, 16'h0000,
16'h21FA, 16'h0000,
16'h21FB, 16'h0000,
16'h21FC, 16'h0000,
16'h21FD, 16'h0000,
16'h21FE, 16'h0000,
16'h21FF, 16'h0000,
16'h2200, 16'h0000,
16'h2201, 16'h0000,
16'h2202, 16'h0000,
16'h2203, 16'h0000,
16'h2204, 16'h0000,
16'h2205, 16'h0000,
16'h2206, 16'h0000,
16'h2207, 16'h0000,
16'h2208, 16'h0000,
16'h2209, 16'h0000,
16'h220A, 16'h0000,
16'h220B, 16'h0000,
16'h220C, 16'h0000,
16'h220D, 16'h0000,
16'h220E, 16'h0000,
16'h220F, 16'h0000,
16'h2210, 16'h0000,
16'h2211, 16'h0000,
16'h2212, 16'h0000,
16'h2213, 16'h0000,
16'h2214, 16'h0000,
16'h2215, 16'h0000,
16'h2216, 16'h0000,
16'h2217, 16'h0000,
16'h2218, 16'h0000,
16'h2219, 16'h0000,
16'h221A, 16'h0000,
16'h221B, 16'h0000,
16'h221C, 16'h0000,
16'h221D, 16'h0000,
16'h221E, 16'h0000,
16'h221F, 16'h0000,
16'h2220, 16'h0000,
16'h2221, 16'h0000,
16'h2222, 16'h0000,
16'h2223, 16'h0000,
16'h2224, 16'h0000,
16'h2225, 16'h0000,
16'h2226, 16'h0000,
16'h2227, 16'h0000,
16'h2228, 16'h0000,
16'h2229, 16'h0000,
16'h222A, 16'h0000,
16'h222B, 16'h0000,
16'h222C, 16'h0000,
16'h222D, 16'h0000,
16'h222E, 16'h0000,
16'h222F, 16'h0000,
16'h2230, 16'h0000,
16'h2231, 16'h0000,
16'h2232, 16'h0000,
16'h2233, 16'h0000,
16'h2234, 16'h0000,
16'h2235, 16'h0000,
16'h2236, 16'h0000,
16'h2237, 16'h0000,
16'h2238, 16'h0000,
16'h2239, 16'h0000,
16'h223A, 16'h0000,
16'h223B, 16'h0000,
16'h223C, 16'h0000,
16'h223D, 16'h0000,
16'h223E, 16'h0000,
16'h223F, 16'h0000,
16'h2240, 16'h0000,
16'h2241, 16'h0000,
16'h2242, 16'h0000,
16'h2243, 16'h0000,
16'h2244, 16'h0000,
16'h2245, 16'h0000,
16'h2246, 16'h0000,
16'h2247, 16'h0000,
16'h2248, 16'h0000,
16'h2249, 16'h0000,
16'h224A, 16'h0000,
16'h224B, 16'h0000,
16'h224C, 16'h0000,
16'h224D, 16'h0000,
16'h224E, 16'h0000,
16'h224F, 16'h0000,
16'h2250, 16'h0000,
16'h2251, 16'h0000,
16'h2252, 16'h0000,
16'h2253, 16'h0000,
16'h2254, 16'h0000,
16'h2255, 16'h0000,
16'h2256, 16'h0000,
16'h2257, 16'h0000,
16'h2258, 16'h0000,
16'h2259, 16'h0000,
16'h225A, 16'h0000,
16'h225B, 16'h0000,
16'h225C, 16'h0000,
16'h225D, 16'h0000,
16'h225E, 16'h0000,
16'h225F, 16'h0000,
16'h2260, 16'h0000,
16'h2261, 16'h0000,
16'h2262, 16'h0000,
16'h2263, 16'h0000,
16'h2264, 16'h0000,
16'h2265, 16'h0000,
16'h2266, 16'h0000,
16'h2267, 16'h0000,
16'h2268, 16'h0000,
16'h2269, 16'h0000,
16'h226A, 16'h0000,
16'h226B, 16'h0000,
16'h226C, 16'h0000,
16'h226D, 16'h0000,
16'h226E, 16'h0000,
16'h226F, 16'h0000,
16'h2270, 16'h0000,
16'h2271, 16'h0000,
16'h2272, 16'h0000,
16'h2273, 16'h0000,
16'h2274, 16'h0000,
16'h2275, 16'h0000,
16'h2276, 16'h0000,
16'h2277, 16'h0000,
16'h2278, 16'h0000,
16'h2279, 16'h0000,
16'h227A, 16'h0000,
16'h227B, 16'h0000,
16'h227C, 16'h0000,
16'h227D, 16'h0000,
16'h227E, 16'h0000,
16'h227F, 16'h0000,
16'h2280, 16'h0000,
16'h2281, 16'h0000,
16'h2282, 16'h0000,
16'h2283, 16'h0000,
16'h2284, 16'h0000,
16'h2285, 16'h0000,
16'h2286, 16'h0000,
16'h2287, 16'h0000,
16'h2288, 16'h0000,
16'h2289, 16'h0000,
16'h228A, 16'h0000,
16'h228B, 16'h0000,
16'h228C, 16'h0000,
16'h228D, 16'h0000,
16'h228E, 16'h0000,
16'h228F, 16'h0000,
16'h2290, 16'h0000,
16'h2291, 16'h0000,
16'h2292, 16'h0000,
16'h2293, 16'h0000,
16'h2294, 16'h0000,
16'h2295, 16'h0000,
16'h2296, 16'h0000,
16'h2297, 16'h0000,
16'h2298, 16'h0000,
16'h2299, 16'h0000,
16'h229A, 16'h0000,
16'h229B, 16'h0000,
16'h229C, 16'h0000,
16'h229D, 16'h0000,
16'h229E, 16'h0000,
16'h229F, 16'h0000,
16'h22A0, 16'h0000,
16'h22A1, 16'h0000,
16'h22A2, 16'h0000,
16'h22A3, 16'h0000,
16'h22A4, 16'h0000,
16'h22A5, 16'h0000,
16'h22A6, 16'h0000,
16'h22A7, 16'h0000,
16'h22A8, 16'h0000,
16'h22A9, 16'h0000,
16'h22AA, 16'h0000,
16'h22AB, 16'h0000,
16'h22AC, 16'h0000,
16'h22AD, 16'h0000,
16'h22AE, 16'h0000,
16'h22AF, 16'h0000,
16'h22B0, 16'h0000,
16'h22B1, 16'h0000,
16'h22B2, 16'h0000,
16'h22B3, 16'h0000,
16'h22B4, 16'h0000,
16'h22B5, 16'h0000,
16'h22B6, 16'h0000,
16'h22B7, 16'h0000,
16'h22B8, 16'h0000,
16'h22B9, 16'h0000,
16'h22BA, 16'h0000,
16'h22BB, 16'h0000,
16'h22BC, 16'h0000,
16'h22BD, 16'h0000,
16'h22BE, 16'h0000,
16'h22BF, 16'h0000,
16'h22C0, 16'h0000,
16'h22C1, 16'h0000,
16'h22C2, 16'h0000,
16'h22C3, 16'h0000,
16'h22C4, 16'h0000,
16'h22C5, 16'h0000,
16'h22C6, 16'h0000,
16'h22C7, 16'h0000,
16'h22C8, 16'h0000,
16'h22C9, 16'h0000,
16'h22CA, 16'h0000,
16'h22CB, 16'h0000,
16'h22CC, 16'h0000,
16'h22CD, 16'h0000,
16'h22CE, 16'h0000,
16'h22CF, 16'h0000,
16'h22D0, 16'h0000,
16'h22D1, 16'h0000,
16'h22D2, 16'h0000,
16'h22D3, 16'h0000,
16'h22D4, 16'h0000,
16'h22D5, 16'h0000,
16'h22D6, 16'h0000,
16'h22D7, 16'h0000,
16'h22D8, 16'h0000,
16'h22D9, 16'h0000,
16'h22DA, 16'h0000,
16'h22DB, 16'h0000,
16'h22DC, 16'h0000,
16'h22DD, 16'h0000,
16'h22DE, 16'h0000,
16'h22DF, 16'h0000,
16'h22E0, 16'h0000,
16'h22E1, 16'h0000,
16'h22E2, 16'h0000,
16'h22E3, 16'h0000,
16'h22E4, 16'h0000,
16'h22E5, 16'h0000,
16'h22E6, 16'h0000,
16'h22E7, 16'h0000,
16'h22E8, 16'h0000,
16'h22E9, 16'h0000,
16'h22EA, 16'h0000,
16'h22EB, 16'h0000,
16'h22EC, 16'h0000,
16'h22ED, 16'h0000,
16'h22EE, 16'h0000,
16'h22EF, 16'h0000,
16'h22F0, 16'h0000,
16'h22F1, 16'h0000,
16'h22F2, 16'h0000,
16'h22F3, 16'h0000,
16'h22F4, 16'h0000,
16'h22F5, 16'h0000,
16'h22F6, 16'h0000,
16'h22F7, 16'h0000,
16'h22F8, 16'h0000,
16'h22F9, 16'h0000,
16'h22FA, 16'h0000,
16'h22FB, 16'h0000,
16'h22FC, 16'h0000,
16'h22FD, 16'h0000,
16'h22FE, 16'h0000,
16'h22FF, 16'h0000,
16'h2300, 16'h0000,
16'h2301, 16'h0000,
16'h2302, 16'h0000,
16'h2303, 16'h0000,
16'h2304, 16'h0000,
16'h2305, 16'h0000,
16'h2306, 16'h0000,
16'h2307, 16'h0000,
16'h2308, 16'h0000,
16'h2309, 16'h0000,
16'h230A, 16'h0000,
16'h230B, 16'h0000,
16'h230C, 16'h0000,
16'h230D, 16'h0000,
16'h230E, 16'h0000,
16'h230F, 16'h0000,
16'h2310, 16'h0000,
16'h2311, 16'h0000,
16'h2312, 16'h0000,
16'h2313, 16'h0000,
16'h2314, 16'h0000,
16'h2315, 16'h0000,
16'h2316, 16'h0000,
16'h2317, 16'h0000,
16'h2318, 16'h0000,
16'h2319, 16'h0000,
16'h231A, 16'h0000,
16'h231B, 16'h0000,
16'h231C, 16'h0000,
16'h231D, 16'h0000,
16'h231E, 16'h0000,
16'h231F, 16'h0000,
16'h2320, 16'h0000,
16'h2321, 16'h0000,
16'h2322, 16'h0000,
16'h2323, 16'h0000,
16'h2324, 16'h0000,
16'h2325, 16'h0000,
16'h2326, 16'h0000,
16'h2327, 16'h0000,
16'h2328, 16'h0000,
16'h2329, 16'h0000,
16'h232A, 16'h0000,
16'h232B, 16'h0000,
16'h232C, 16'h0000,
16'h232D, 16'h0000,
16'h232E, 16'h0000,
16'h232F, 16'h0000,
16'h2330, 16'h0000,
16'h2331, 16'h0000,
16'h2332, 16'h0000,
16'h2333, 16'h0000,
16'h2334, 16'h0000,
16'h2335, 16'h0000,
16'h2336, 16'h0000,
16'h2337, 16'h0000,
16'h2338, 16'h0000,
16'h2339, 16'h0000,
16'h233A, 16'h0000,
16'h233B, 16'h0000,
16'h233C, 16'h0000,
16'h233D, 16'h0000,
16'h233E, 16'h0000,
16'h233F, 16'h0000,
16'h2340, 16'h0000,
16'h2341, 16'h0000,
16'h2342, 16'h0000,
16'h2343, 16'h0000,
16'h2344, 16'h0000,
16'h2345, 16'h0000,
16'h2346, 16'h0000,
16'h2347, 16'h0000,
16'h2348, 16'h0000,
16'h2349, 16'h0000,
16'h234A, 16'h0000,
16'h234B, 16'h0000,
16'h234C, 16'h0000,
16'h234D, 16'h0000,
16'h234E, 16'h0000,
16'h234F, 16'h0000,
16'h2350, 16'h0000,
16'h2351, 16'h0000,
16'h2352, 16'h0000,
16'h2353, 16'h0000,
16'h2354, 16'h0000,
16'h2355, 16'h0000,
16'h2356, 16'h0000,
16'h2357, 16'h0000,
16'h2358, 16'h0000,
16'h2359, 16'h0000,
16'h235A, 16'h0000,
16'h235B, 16'h0000,
16'h235C, 16'h0000,
16'h235D, 16'h0000,
16'h235E, 16'h0000,
16'h235F, 16'h0000,
16'h2360, 16'h0000,
16'h2361, 16'h0000,
16'h2362, 16'h0000,
16'h2363, 16'h0000,
16'h2364, 16'h0000,
16'h2365, 16'h0000,
16'h2366, 16'h0000,
16'h2367, 16'h0000,
16'h2368, 16'h0000,
16'h2369, 16'h0000,
16'h236A, 16'h0000,
16'h236B, 16'h0000,
16'h236C, 16'h0000,
16'h236D, 16'h0000,
16'h236E, 16'h0000,
16'h236F, 16'h0000,
16'h2370, 16'h0000,
16'h2371, 16'h0000,
16'h2372, 16'h0000,
16'h2373, 16'h0000,
16'h2374, 16'h0000,
16'h2375, 16'h0000,
16'h2376, 16'h0000,
16'h2377, 16'h0000,
16'h2378, 16'h0000,
16'h2379, 16'h0000,
16'h237A, 16'h0000,
16'h237B, 16'h0000,
16'h237C, 16'h0000,
16'h237D, 16'h0000,
16'h237E, 16'h0000,
16'h237F, 16'h0000,
16'h2380, 16'h0000,
16'h2381, 16'h0000,
16'h2382, 16'h0000,
16'h2383, 16'h0000,
16'h2384, 16'h0000,
16'h2385, 16'h0000,
16'h2386, 16'h0000,
16'h2387, 16'h0000,
16'h2388, 16'h0000,
16'h2389, 16'h0000,
16'h238A, 16'h0000,
16'h238B, 16'h0000,
16'h238C, 16'h0000,
16'h238D, 16'h0000,
16'h238E, 16'h0000,
16'h238F, 16'h0000,
16'h2390, 16'h0000,
16'h2391, 16'h0000,
16'h2392, 16'h0000,
16'h2393, 16'h0000,
16'h2394, 16'h0000,
16'h2395, 16'h0000,
16'h2396, 16'h0000,
16'h2397, 16'h0000,
16'h2398, 16'h0000,
16'h2399, 16'h0000,
16'h239A, 16'h0000,
16'h239B, 16'h0000,
16'h239C, 16'h0000,
16'h239D, 16'h0000,
16'h239E, 16'h0000,
16'h239F, 16'h0000,
16'h23A0, 16'h0000,
16'h23A1, 16'h0000,
16'h23A2, 16'h0000,
16'h23A3, 16'h0000,
16'h23A4, 16'h0000,
16'h23A5, 16'h0000,
16'h23A6, 16'h0000,
16'h23A7, 16'h0000,
16'h23A8, 16'h0000,
16'h23A9, 16'h0000,
16'h23AA, 16'h0000,
16'h23AB, 16'h0000,
16'h23AC, 16'h0000,
16'h23AD, 16'h0000,
16'h23AE, 16'h0000,
16'h23AF, 16'h0000,
16'h23B0, 16'h0000,
16'h23B1, 16'h0000,
16'h23B2, 16'h0000,
16'h23B3, 16'h0000,
16'h23B4, 16'h0000,
16'h23B5, 16'h0000,
16'h23B6, 16'h0000,
16'h23B7, 16'h0000,
16'h23B8, 16'h0000,
16'h23B9, 16'h0000,
16'h23BA, 16'h0000,
16'h23BB, 16'h0000,
16'h23BC, 16'h0000,
16'h23BD, 16'h0000,
16'h23BE, 16'h0000,
16'h23BF, 16'h0000,
16'h23C0, 16'h0000,
16'h23C1, 16'h0000,
16'h23C2, 16'h0000,
16'h23C3, 16'h0000,
16'h23C4, 16'h0000,
16'h23C5, 16'h0000,
16'h23C6, 16'h0000,
16'h23C7, 16'h0000,
16'h23C8, 16'h0000,
16'h23C9, 16'h0000,
16'h23CA, 16'h0000,
16'h23CB, 16'h0000,
16'h23CC, 16'h0000,
16'h23CD, 16'h0000,
16'h23CE, 16'h0000,
16'h23CF, 16'h0000,
16'h23D0, 16'h0000,
16'h23D1, 16'h0000,
16'h23D2, 16'h0000,
16'h23D3, 16'h0000,
16'h23D4, 16'h0000,
16'h23D5, 16'h0000,
16'h23D6, 16'h0000,
16'h23D7, 16'h0000,
16'h23D8, 16'h0000,
16'h23D9, 16'h0000,
16'h23DA, 16'h0000,
16'h23DB, 16'h0000,
16'h23DC, 16'h0000,
16'h23DD, 16'h0000,
16'h23DE, 16'h0000,
16'h23DF, 16'h0000,
16'h23E0, 16'h0000,
16'h23E1, 16'h0000,
16'h23E2, 16'h0000,
16'h23E3, 16'h0000,
16'h23E4, 16'h0000,
16'h23E5, 16'h0000,
16'h23E6, 16'h0000,
16'h23E7, 16'h0000,
16'h23E8, 16'h0000,
16'h23E9, 16'h0000,
16'h23EA, 16'h0000,
16'h23EB, 16'h0000,
16'h23EC, 16'h0000,
16'h23ED, 16'h0000,
16'h23EE, 16'h0000,
16'h23EF, 16'h0000,
16'h23F0, 16'h0000,
16'h23F1, 16'h0000,
16'h23F2, 16'h0000,
16'h23F3, 16'h0000,
16'h23F4, 16'h0000,
16'h23F5, 16'h0000,
16'h23F6, 16'h0000,
16'h23F7, 16'h0000,
16'h23F8, 16'h0000,
16'h23F9, 16'h0000,
16'h23FA, 16'h0000,
16'h23FB, 16'h0000,
16'h23FC, 16'h0000,
16'h23FD, 16'h0000,
16'h23FE, 16'h0000,
16'h23FF, 16'h0000,
16'h2400, 16'h0001,
16'h2401, 16'h0001,
16'h2402, 16'h0001,
16'h2403, 16'h0001,
16'h2404, 16'h0001,
16'h2405, 16'h0001,
16'h2406, 16'h0001,
16'h2407, 16'h0001,
16'h2408, 16'h0001,
16'h2409, 16'h0001,
16'h240A, 16'h0001,
16'h240B, 16'h0001,
16'h240C, 16'h0001,
16'h240D, 16'h0001,
16'h240E, 16'h0001,
16'h240F, 16'h0001,
16'h2410, 16'h0001,
16'h2411, 16'h0001,
16'h2412, 16'h0001,
16'h2413, 16'h0001,
16'h2414, 16'h0001,
16'h2415, 16'h0001,
16'h2416, 16'h0001,
16'h2417, 16'h0001,
16'h2418, 16'h0001,
16'h2419, 16'h0001,
16'h241A, 16'h0001,
16'h241B, 16'h0001,
16'h241C, 16'h0001,
16'h241D, 16'h0001,
16'h241E, 16'h0001,
16'h241F, 16'h0001,
16'h2420, 16'h0001,
16'h2421, 16'h0001,
16'h2422, 16'h0001,
16'h2423, 16'h0001,
16'h2424, 16'h0001,
16'h2425, 16'h0001,
16'h2426, 16'h0001,
16'h2427, 16'h0001,
16'h2428, 16'h0001,
16'h2429, 16'h0001,
16'h242A, 16'h0001,
16'h242B, 16'h0001,
16'h242C, 16'h0001,
16'h242D, 16'h0001,
16'h242E, 16'h0001,
16'h242F, 16'h0001,
16'h2430, 16'h0001,
16'h2431, 16'h0001,
16'h2432, 16'h0001,
16'h2433, 16'h0001,
16'h2434, 16'h0001,
16'h2435, 16'h0001,
16'h2436, 16'h0001,
16'h2437, 16'h0001,
16'h2438, 16'h0001,
16'h2439, 16'h0001,
16'h243A, 16'h0001,
16'h243B, 16'h0001,
16'h243C, 16'h0001,
16'h243D, 16'h0001,
16'h243E, 16'h0001,
16'h243F, 16'h0001,
16'h2440, 16'h0001,
16'h2441, 16'h0001,
16'h2442, 16'h0001,
16'h2443, 16'h0001,
16'h2444, 16'h0001,
16'h2445, 16'h0001,
16'h2446, 16'h0001,
16'h2447, 16'h0001,
16'h2448, 16'h0001,
16'h2449, 16'h0001,
16'h244A, 16'h0001,
16'h244B, 16'h0001,
16'h244C, 16'h0001,
16'h244D, 16'h0001,
16'h244E, 16'h0001,
16'h244F, 16'h0001,
16'h2450, 16'h0001,
16'h2451, 16'h0001,
16'h2452, 16'h0001,
16'h2453, 16'h0001,
16'h2454, 16'h0001,
16'h2455, 16'h0001,
16'h2456, 16'h0001,
16'h2457, 16'h0001,
16'h2458, 16'h0001,
16'h2459, 16'h0001,
16'h245A, 16'h0001,
16'h245B, 16'h0001,
16'h245C, 16'h0001,
16'h245D, 16'h0001,
16'h245E, 16'h0001,
16'h245F, 16'h0001,
16'h2460, 16'h0001,
16'h2461, 16'h0001,
16'h2462, 16'h0001,
16'h2463, 16'h0001,
16'h2464, 16'h0001,
16'h2465, 16'h0001,
16'h2466, 16'h0001,
16'h2467, 16'h0001,
16'h2468, 16'h0001,
16'h2469, 16'h0001,
16'h246A, 16'h0001,
16'h246B, 16'h0001,
16'h246C, 16'h0001,
16'h246D, 16'h0001,
16'h246E, 16'h0001,
16'h246F, 16'h0001,
16'h2470, 16'h0001,
16'h2471, 16'h0001,
16'h2472, 16'h0001,
16'h2473, 16'h0001,
16'h2474, 16'h0001,
16'h2475, 16'h0001,
16'h2476, 16'h0001,
16'h2477, 16'h0001,
16'h2478, 16'h0001,
16'h2479, 16'h0001,
16'h247A, 16'h0001,
16'h247B, 16'h0001,
16'h247C, 16'h0001,
16'h247D, 16'h0001,
16'h247E, 16'h0001,
16'h247F, 16'h0001,
16'h2480, 16'h0001,
16'h2481, 16'h0001,
16'h2482, 16'h0001,
16'h2483, 16'h0001,
16'h2484, 16'h0001,
16'h2485, 16'h0001,
16'h2486, 16'h0001,
16'h2487, 16'h0001,
16'h2488, 16'h0001,
16'h2489, 16'h0001,
16'h248A, 16'h0001,
16'h248B, 16'h0001,
16'h248C, 16'h0001,
16'h248D, 16'h0001,
16'h248E, 16'h0001,
16'h248F, 16'h0001,
16'h2490, 16'h0001,
16'h2491, 16'h0001,
16'h2492, 16'h0001,
16'h2493, 16'h0001,
16'h2494, 16'h0001,
16'h2495, 16'h0001,
16'h2496, 16'h0001,
16'h2497, 16'h0001,
16'h2498, 16'h0001,
16'h2499, 16'h0001,
16'h249A, 16'h0001,
16'h249B, 16'h0001,
16'h249C, 16'h0001,
16'h249D, 16'h0001,
16'h249E, 16'h0001,
16'h249F, 16'h0001,
16'h24A0, 16'h0001,
16'h24A1, 16'h0001,
16'h24A2, 16'h0001,
16'h24A3, 16'h0001,
16'h24A4, 16'h0001,
16'h24A5, 16'h0001,
16'h24A6, 16'h0001,
16'h24A7, 16'h0001,
16'h24A8, 16'h0001,
16'h24A9, 16'h0001,
16'h24AA, 16'h0001,
16'h24AB, 16'h0001,
16'h24AC, 16'h0001,
16'h24AD, 16'h0001,
16'h24AE, 16'h0001,
16'h24AF, 16'h0001,
16'h24B0, 16'h0001,
16'h24B1, 16'h0001,
16'h24B2, 16'h0001,
16'h24B3, 16'h0001,
16'h24B4, 16'h0001,
16'h24B5, 16'h0001,
16'h24B6, 16'h0001,
16'h24B7, 16'h0001,
16'h24B8, 16'h0001,
16'h24B9, 16'h0001,
16'h24BA, 16'h0001,
16'h24BB, 16'h0001,
16'h24BC, 16'h0001,
16'h24BD, 16'h0001,
16'h24BE, 16'h0001,
16'h24BF, 16'h0001,
16'h24C0, 16'h0001,
16'h24C1, 16'h0001,
16'h24C2, 16'h0001,
16'h24C3, 16'h0001,
16'h24C4, 16'h0001,
16'h24C5, 16'h0001,
16'h24C6, 16'h0001,
16'h24C7, 16'h0001,
16'h24C8, 16'h0001,
16'h24C9, 16'h0001,
16'h24CA, 16'h0001,
16'h24CB, 16'h0001,
16'h24CC, 16'h0001,
16'h24CD, 16'h0001,
16'h24CE, 16'h0001,
16'h24CF, 16'h0001,
16'h24D0, 16'h0001,
16'h24D1, 16'h0001,
16'h24D2, 16'h0001,
16'h24D3, 16'h0001,
16'h24D4, 16'h0001,
16'h24D5, 16'h0001,
16'h24D6, 16'h0001,
16'h24D7, 16'h0001,
16'h24D8, 16'h0001,
16'h24D9, 16'h0001,
16'h24DA, 16'h0001,
16'h24DB, 16'h0001,
16'h24DC, 16'h0001,
16'h24DD, 16'h0001,
16'h24DE, 16'h0001,
16'h24DF, 16'h0001,
16'h24E0, 16'h0001,
16'h24E1, 16'h0001,
16'h24E2, 16'h0001,
16'h24E3, 16'h0001,
16'h24E4, 16'h0001,
16'h24E5, 16'h0001,
16'h24E6, 16'h0001,
16'h24E7, 16'h0001,
16'h24E8, 16'h0001,
16'h24E9, 16'h0001,
16'h24EA, 16'h0001,
16'h24EB, 16'h0001,
16'h24EC, 16'h0001,
16'h24ED, 16'h0001,
16'h24EE, 16'h0001,
16'h24EF, 16'h0001,
16'h24F0, 16'h0001,
16'h24F1, 16'h0001,
16'h24F2, 16'h0001,
16'h24F3, 16'h0001,
16'h24F4, 16'h0001,
16'h24F5, 16'h0001,
16'h24F6, 16'h0001,
16'h24F7, 16'h0001,
16'h24F8, 16'h0001,
16'h24F9, 16'h0001,
16'h24FA, 16'h0001,
16'h24FB, 16'h0001,
16'h24FC, 16'h0001,
16'h24FD, 16'h0001,
16'h24FE, 16'h0001,
16'h24FF, 16'h0001,
16'h2500, 16'h0001,
16'h2501, 16'h0001,
16'h2502, 16'h0001,
16'h2503, 16'h0001,
16'h2504, 16'h0001,
16'h2505, 16'h0001,
16'h2506, 16'h0001,
16'h2507, 16'h0001,
16'h2508, 16'h0001,
16'h2509, 16'h0001,
16'h250A, 16'h0001,
16'h250B, 16'h0001,
16'h250C, 16'h0001,
16'h250D, 16'h0001,
16'h250E, 16'h0001,
16'h250F, 16'h0001,
16'h2510, 16'h0001,
16'h2511, 16'h0001,
16'h2512, 16'h0001,
16'h2513, 16'h0001,
16'h2514, 16'h0001,
16'h2515, 16'h0001,
16'h2516, 16'h0001,
16'h2517, 16'h0001,
16'h2518, 16'h0001,
16'h2519, 16'h0001,
16'h251A, 16'h0001,
16'h251B, 16'h0001,
16'h251C, 16'h0001,
16'h251D, 16'h0001,
16'h251E, 16'h0001,
16'h251F, 16'h0001,
16'h2520, 16'h0001,
16'h2521, 16'h0001,
16'h2522, 16'h0001,
16'h2523, 16'h0001,
16'h2524, 16'h0001,
16'h2525, 16'h0001,
16'h2526, 16'h0001,
16'h2527, 16'h0001,
16'h2528, 16'h0001,
16'h2529, 16'h0001,
16'h252A, 16'h0001,
16'h252B, 16'h0001,
16'h252C, 16'h0001,
16'h252D, 16'h0001,
16'h252E, 16'h0001,
16'h252F, 16'h0001,
16'h2530, 16'h0001,
16'h2531, 16'h0001,
16'h2532, 16'h0001,
16'h2533, 16'h0001,
16'h2534, 16'h0001,
16'h2535, 16'h0001,
16'h2536, 16'h0001,
16'h2537, 16'h0001,
16'h2538, 16'h0001,
16'h2539, 16'h0001,
16'h253A, 16'h0001,
16'h253B, 16'h0001,
16'h253C, 16'h0001,
16'h253D, 16'h0001,
16'h253E, 16'h0001,
16'h253F, 16'h0001,
16'h2540, 16'h0001,
16'h2541, 16'h0001,
16'h2542, 16'h0001,
16'h2543, 16'h0001,
16'h2544, 16'h0001,
16'h2545, 16'h0001,
16'h2546, 16'h0001,
16'h2547, 16'h0001,
16'h2548, 16'h0001,
16'h2549, 16'h0001,
16'h254A, 16'h0001,
16'h254B, 16'h0001,
16'h254C, 16'h0001,
16'h254D, 16'h0001,
16'h254E, 16'h0001,
16'h254F, 16'h0001,
16'h2550, 16'h0001,
16'h2551, 16'h0001,
16'h2552, 16'h0001,
16'h2553, 16'h0001,
16'h2554, 16'h0001,
16'h2555, 16'h0001,
16'h2556, 16'h0001,
16'h2557, 16'h0001,
16'h2558, 16'h0001,
16'h2559, 16'h0001,
16'h255A, 16'h0001,
16'h255B, 16'h0001,
16'h255C, 16'h0001,
16'h255D, 16'h0001,
16'h255E, 16'h0001,
16'h255F, 16'h0001,
16'h2560, 16'h0001,
16'h2561, 16'h0001,
16'h2562, 16'h0001,
16'h2563, 16'h0001,
16'h2564, 16'h0001,
16'h2565, 16'h0001,
16'h2566, 16'h0001,
16'h2567, 16'h0001,
16'h2568, 16'h0001,
16'h2569, 16'h0001,
16'h256A, 16'h0001,
16'h256B, 16'h0001,
16'h256C, 16'h0001,
16'h256D, 16'h0001,
16'h256E, 16'h0001,
16'h256F, 16'h0001,
16'h2570, 16'h0001,
16'h2571, 16'h0001,
16'h2572, 16'h0001,
16'h2573, 16'h0001,
16'h2574, 16'h0001,
16'h2575, 16'h0001,
16'h2576, 16'h0001,
16'h2577, 16'h0001,
16'h2578, 16'h0001,
16'h2579, 16'h0001,
16'h257A, 16'h0001,
16'h257B, 16'h0001,
16'h257C, 16'h0001,
16'h257D, 16'h0001,
16'h257E, 16'h0001,
16'h257F, 16'h0001,
16'h2580, 16'h0001,
16'h2581, 16'h0001,
16'h2582, 16'h0001,
16'h2583, 16'h0001,
16'h2584, 16'h0001,
16'h2585, 16'h0001,
16'h2586, 16'h0001,
16'h2587, 16'h0001,
16'h2588, 16'h0001,
16'h2589, 16'h0001,
16'h258A, 16'h0001,
16'h258B, 16'h0001,
16'h258C, 16'h0001,
16'h258D, 16'h0001,
16'h258E, 16'h0001,
16'h258F, 16'h0001,
16'h2590, 16'h0001,
16'h2591, 16'h0001,
16'h2592, 16'h0001,
16'h2593, 16'h0001,
16'h2594, 16'h0001,
16'h2595, 16'h0001,
16'h2596, 16'h0001,
16'h2597, 16'h0001,
16'h2598, 16'h0001,
16'h2599, 16'h0001,
16'h259A, 16'h0001,
16'h259B, 16'h0001,
16'h259C, 16'h0001,
16'h259D, 16'h0001,
16'h259E, 16'h0001,
16'h259F, 16'h0001,
16'h25A0, 16'h0001,
16'h25A1, 16'h0001,
16'h25A2, 16'h0001,
16'h25A3, 16'h0001,
16'h25A4, 16'h0001,
16'h25A5, 16'h0001,
16'h25A6, 16'h0001,
16'h25A7, 16'h0001,
16'h25A8, 16'h0001,
16'h25A9, 16'h0001,
16'h25AA, 16'h0001,
16'h25AB, 16'h0001,
16'h25AC, 16'h0001,
16'h25AD, 16'h0001,
16'h25AE, 16'h0001,
16'h25AF, 16'h0001,
16'h25B0, 16'h0001,
16'h25B1, 16'h0001,
16'h25B2, 16'h0001,
16'h25B3, 16'h0001,
16'h25B4, 16'h0001,
16'h25B5, 16'h0001,
16'h25B6, 16'h0001,
16'h25B7, 16'h0001,
16'h25B8, 16'h0001,
16'h25B9, 16'h0001,
16'h25BA, 16'h0001,
16'h25BB, 16'h0001,
16'h25BC, 16'h0001,
16'h25BD, 16'h0001,
16'h25BE, 16'h0001,
16'h25BF, 16'h0001,
16'h25C0, 16'h0001,
16'h25C1, 16'h0001,
16'h25C2, 16'h0001,
16'h25C3, 16'h0001,
16'h25C4, 16'h0001,
16'h25C5, 16'h0001,
16'h25C6, 16'h0001,
16'h25C7, 16'h0001,
16'h25C8, 16'h0001,
16'h25C9, 16'h0001,
16'h25CA, 16'h0001,
16'h25CB, 16'h0001,
16'h25CC, 16'h0001,
16'h25CD, 16'h0001,
16'h25CE, 16'h0001,
16'h25CF, 16'h0001,
16'h25D0, 16'h0001,
16'h25D1, 16'h0001,
16'h25D2, 16'h0001,
16'h25D3, 16'h0001,
16'h25D4, 16'h0001,
16'h25D5, 16'h0001,
16'h25D6, 16'h0001,
16'h25D7, 16'h0001,
16'h25D8, 16'h0001,
16'h25D9, 16'h0001,
16'h25DA, 16'h0001,
16'h25DB, 16'h0001,
16'h25DC, 16'h0001,
16'h25DD, 16'h0001,
16'h25DE, 16'h0001,
16'h25DF, 16'h0001,
16'h25E0, 16'h0001,
16'h25E1, 16'h0001,
16'h25E2, 16'h0001,
16'h25E3, 16'h0001,
16'h25E4, 16'h0001,
16'h25E5, 16'h0001,
16'h25E6, 16'h0001,
16'h25E7, 16'h0001,
16'h25E8, 16'h0001,
16'h25E9, 16'h0001,
16'h25EA, 16'h0001,
16'h25EB, 16'h0001,
16'h25EC, 16'h0001,
16'h25ED, 16'h0001,
16'h25EE, 16'h0001,
16'h25EF, 16'h0001,
16'h25F0, 16'h0001,
16'h25F1, 16'h0001,
16'h25F2, 16'h0001,
16'h25F3, 16'h0001,
16'h25F4, 16'h0001,
16'h25F5, 16'h0001,
16'h25F6, 16'h0001,
16'h25F7, 16'h0001,
16'h25F8, 16'h0001,
16'h25F9, 16'h0001,
16'h25FA, 16'h0001,
16'h25FB, 16'h0001,
16'h25FC, 16'h0001,
16'h25FD, 16'h0001,
16'h25FE, 16'h0001,
16'h25FF, 16'h0001,
16'h2600, 16'h0001,
16'h2601, 16'h0001,
16'h2602, 16'h0001,
16'h2603, 16'h0001,
16'h2604, 16'h0001,
16'h2605, 16'h0001,
16'h2606, 16'h0001,
16'h2607, 16'h0001,
16'h2608, 16'h0001,
16'h2609, 16'h0001,
16'h260A, 16'h0001,
16'h260B, 16'h0001,
16'h260C, 16'h0001,
16'h260D, 16'h0001,
16'h260E, 16'h0001,
16'h260F, 16'h0001,
16'h2610, 16'h0001,
16'h2611, 16'h0001,
16'h2612, 16'h0001,
16'h2613, 16'h0001,
16'h2614, 16'h0001,
16'h2615, 16'h0001,
16'h2616, 16'h0001,
16'h2617, 16'h0001,
16'h2618, 16'h0001,
16'h2619, 16'h0001,
16'h261A, 16'h0001,
16'h261B, 16'h0001,
16'h261C, 16'h0001,
16'h261D, 16'h0001,
16'h261E, 16'h0001,
16'h261F, 16'h0001,
16'h2620, 16'h0001,
16'h2621, 16'h0001,
16'h2622, 16'h0001,
16'h2623, 16'h0001,
16'h2624, 16'h0001,
16'h2625, 16'h0001,
16'h2626, 16'h0001,
16'h2627, 16'h0001,
16'h2628, 16'h0001,
16'h2629, 16'h0001,
16'h262A, 16'h0001,
16'h262B, 16'h0001,
16'h262C, 16'h0001,
16'h262D, 16'h0001,
16'h262E, 16'h0001,
16'h262F, 16'h0001,
16'h2630, 16'h0001,
16'h2631, 16'h0001,
16'h2632, 16'h0001,
16'h2633, 16'h0001,
16'h2634, 16'h0001,
16'h2635, 16'h0001,
16'h2636, 16'h0001,
16'h2637, 16'h0001,
16'h2638, 16'h0001,
16'h2639, 16'h0001,
16'h263A, 16'h0001,
16'h263B, 16'h0001,
16'h263C, 16'h0001,
16'h263D, 16'h0001,
16'h263E, 16'h0001,
16'h263F, 16'h0001,
16'h2640, 16'h0001,
16'h2641, 16'h0001,
16'h2642, 16'h0001,
16'h2643, 16'h0001,
16'h2644, 16'h0001,
16'h2645, 16'h0001,
16'h2646, 16'h0001,
16'h2647, 16'h0001,
16'h2648, 16'h0001,
16'h2649, 16'h0001,
16'h264A, 16'h0001,
16'h264B, 16'h0001,
16'h264C, 16'h0001,
16'h264D, 16'h0001,
16'h264E, 16'h0001,
16'h264F, 16'h0001,
16'h2650, 16'h0001,
16'h2651, 16'h0001,
16'h2652, 16'h0001,
16'h2653, 16'h0001,
16'h2654, 16'h0001,
16'h2655, 16'h0001,
16'h2656, 16'h0001,
16'h2657, 16'h0001,
16'h2658, 16'h0001,
16'h2659, 16'h0001,
16'h265A, 16'h0001,
16'h265B, 16'h0001,
16'h265C, 16'h0001,
16'h265D, 16'h0001,
16'h265E, 16'h0001,
16'h265F, 16'h0001,
16'h2660, 16'h0001,
16'h2661, 16'h0001,
16'h2662, 16'h0001,
16'h2663, 16'h0001,
16'h2664, 16'h0001,
16'h2665, 16'h0001,
16'h2666, 16'h0001,
16'h2667, 16'h0001,
16'h2668, 16'h0001,
16'h2669, 16'h0001,
16'h266A, 16'h0001,
16'h266B, 16'h0001,
16'h266C, 16'h0001,
16'h266D, 16'h0001,
16'h266E, 16'h0001,
16'h266F, 16'h0001,
16'h2670, 16'h0001,
16'h2671, 16'h0001,
16'h2672, 16'h0001,
16'h2673, 16'h0001,
16'h2674, 16'h0001,
16'h2675, 16'h0001,
16'h2676, 16'h0001,
16'h2677, 16'h0001,
16'h2678, 16'h0001,
16'h2679, 16'h0001,
16'h267A, 16'h0001,
16'h267B, 16'h0001,
16'h267C, 16'h0001,
16'h267D, 16'h0001,
16'h267E, 16'h0001,
16'h267F, 16'h0001,
16'h2680, 16'h0001,
16'h2681, 16'h0001,
16'h2682, 16'h0001,
16'h2683, 16'h0001,
16'h2684, 16'h0001,
16'h2685, 16'h0001,
16'h2686, 16'h0001,
16'h2687, 16'h0001,
16'h2688, 16'h0001,
16'h2689, 16'h0001,
16'h268A, 16'h0001,
16'h268B, 16'h0001,
16'h268C, 16'h0001,
16'h268D, 16'h0001,
16'h268E, 16'h0001,
16'h268F, 16'h0001,
16'h2690, 16'h0001,
16'h2691, 16'h0001,
16'h2692, 16'h0001,
16'h2693, 16'h0001,
16'h2694, 16'h0001,
16'h2695, 16'h0001,
16'h2696, 16'h0001,
16'h2697, 16'h0001,
16'h2698, 16'h0001,
16'h2699, 16'h0001,
16'h269A, 16'h0001,
16'h269B, 16'h0001,
16'h269C, 16'h0001,
16'h269D, 16'h0001,
16'h269E, 16'h0001,
16'h269F, 16'h0001,
16'h26A0, 16'h0001,
16'h26A1, 16'h0001,
16'h26A2, 16'h0001,
16'h26A3, 16'h0001,
16'h26A4, 16'h0001,
16'h26A5, 16'h0001,
16'h26A6, 16'h0001,
16'h26A7, 16'h0001,
16'h26A8, 16'h0001,
16'h26A9, 16'h0001,
16'h26AA, 16'h0001,
16'h26AB, 16'h0001,
16'h26AC, 16'h0001,
16'h26AD, 16'h0001,
16'h26AE, 16'h0001,
16'h26AF, 16'h0001,
16'h26B0, 16'h0001,
16'h26B1, 16'h0001,
16'h26B2, 16'h0001,
16'h26B3, 16'h0001,
16'h26B4, 16'h0001,
16'h26B5, 16'h0001,
16'h26B6, 16'h0001,
16'h26B7, 16'h0001,
16'h26B8, 16'h0001,
16'h26B9, 16'h0001,
16'h26BA, 16'h0001,
16'h26BB, 16'h0001,
16'h26BC, 16'h0001,
16'h26BD, 16'h0001,
16'h26BE, 16'h0001,
16'h26BF, 16'h0001,
16'h26C0, 16'h0001,
16'h26C1, 16'h0001,
16'h26C2, 16'h0001,
16'h26C3, 16'h0001,
16'h26C4, 16'h0001,
16'h26C5, 16'h0001,
16'h26C6, 16'h0001,
16'h26C7, 16'h0001,
16'h26C8, 16'h0001,
16'h26C9, 16'h0001,
16'h26CA, 16'h0001,
16'h26CB, 16'h0001,
16'h26CC, 16'h0001,
16'h26CD, 16'h0001,
16'h26CE, 16'h0001,
16'h26CF, 16'h0001,
16'h26D0, 16'h0001,
16'h26D1, 16'h0001,
16'h26D2, 16'h0001,
16'h26D3, 16'h0001,
16'h26D4, 16'h0001,
16'h26D5, 16'h0001,
16'h26D6, 16'h0001,
16'h26D7, 16'h0001,
16'h26D8, 16'h0001,
16'h26D9, 16'h0001,
16'h26DA, 16'h0001,
16'h26DB, 16'h0001,
16'h26DC, 16'h0001,
16'h26DD, 16'h0001,
16'h26DE, 16'h0001,
16'h26DF, 16'h0001,
16'h26E0, 16'h0001,
16'h26E1, 16'h0001,
16'h26E2, 16'h0001,
16'h26E3, 16'h0001,
16'h26E4, 16'h0001,
16'h26E5, 16'h0001,
16'h26E6, 16'h0001,
16'h26E7, 16'h0001,
16'h26E8, 16'h0001,
16'h26E9, 16'h0001,
16'h26EA, 16'h0001,
16'h26EB, 16'h0001,
16'h26EC, 16'h0001,
16'h26ED, 16'h0001,
16'h26EE, 16'h0001,
16'h26EF, 16'h0001,
16'h26F0, 16'h0001,
16'h26F1, 16'h0001,
16'h26F2, 16'h0001,
16'h26F3, 16'h0001,
16'h26F4, 16'h0001,
16'h26F5, 16'h0001,
16'h26F6, 16'h0001,
16'h26F7, 16'h0001,
16'h26F8, 16'h0001,
16'h26F9, 16'h0001,
16'h26FA, 16'h0001,
16'h26FB, 16'h0001,
16'h26FC, 16'h0001,
16'h26FD, 16'h0001,
16'h26FE, 16'h0001,
16'h26FF, 16'h0001,
16'h2700, 16'h0001,
16'h2701, 16'h0001,
16'h2702, 16'h0001,
16'h2703, 16'h0001,
16'h2704, 16'h0001,
16'h2705, 16'h0001,
16'h2706, 16'h0001,
16'h2707, 16'h0001,
16'h2708, 16'h0001,
16'h2709, 16'h0001,
16'h270A, 16'h0001,
16'h270B, 16'h0001,
16'h270C, 16'h0001,
16'h270D, 16'h0001,
16'h270E, 16'h0001,
16'h270F, 16'h0001,
16'h2710, 16'h0001,
16'h2711, 16'h0001,
16'h2712, 16'h0001,
16'h2713, 16'h0001,
16'h2714, 16'h0001,
16'h2715, 16'h0001,
16'h2716, 16'h0001,
16'h2717, 16'h0001,
16'h2718, 16'h0001,
16'h2719, 16'h0001,
16'h271A, 16'h0001,
16'h271B, 16'h0001,
16'h271C, 16'h0001,
16'h271D, 16'h0001,
16'h271E, 16'h0001,
16'h271F, 16'h0001,
16'h2720, 16'h0001,
16'h2721, 16'h0001,
16'h2722, 16'h0001,
16'h2723, 16'h0001,
16'h2724, 16'h0001,
16'h2725, 16'h0001,
16'h2726, 16'h0001,
16'h2727, 16'h0001,
16'h2728, 16'h0001,
16'h2729, 16'h0001,
16'h272A, 16'h0001,
16'h272B, 16'h0001,
16'h272C, 16'h0001,
16'h272D, 16'h0001,
16'h272E, 16'h0001,
16'h272F, 16'h0001,
16'h2730, 16'h0001,
16'h2731, 16'h0001,
16'h2732, 16'h0001,
16'h2733, 16'h0001,
16'h2734, 16'h0001,
16'h2735, 16'h0001,
16'h2736, 16'h0001,
16'h2737, 16'h0001,
16'h2738, 16'h0001,
16'h2739, 16'h0001,
16'h273A, 16'h0001,
16'h273B, 16'h0001,
16'h273C, 16'h0001,
16'h273D, 16'h0001,
16'h273E, 16'h0001,
16'h273F, 16'h0001,
16'h2740, 16'h0001,
16'h2741, 16'h0001,
16'h2742, 16'h0001,
16'h2743, 16'h0001,
16'h2744, 16'h0001,
16'h2745, 16'h0001,
16'h2746, 16'h0001,
16'h2747, 16'h0001,
16'h2748, 16'h0001,
16'h2749, 16'h0001,
16'h274A, 16'h0001,
16'h274B, 16'h0001,
16'h274C, 16'h0001,
16'h274D, 16'h0001,
16'h274E, 16'h0001,
16'h274F, 16'h0001,
16'h2750, 16'h0001,
16'h2751, 16'h0001,
16'h2752, 16'h0001,
16'h2753, 16'h0001,
16'h2754, 16'h0001,
16'h2755, 16'h0001,
16'h2756, 16'h0001,
16'h2757, 16'h0001,
16'h2758, 16'h0001,
16'h2759, 16'h0001,
16'h275A, 16'h0001,
16'h275B, 16'h0001,
16'h275C, 16'h0001,
16'h275D, 16'h0001,
16'h275E, 16'h0001,
16'h275F, 16'h0001,
16'h2760, 16'h0001,
16'h2761, 16'h0001,
16'h2762, 16'h0001,
16'h2763, 16'h0001,
16'h2764, 16'h0001,
16'h2765, 16'h0001,
16'h2766, 16'h0001,
16'h2767, 16'h0001,
16'h2768, 16'h0001,
16'h2769, 16'h0001,
16'h276A, 16'h0001,
16'h276B, 16'h0001,
16'h276C, 16'h0001,
16'h276D, 16'h0001,
16'h276E, 16'h0001,
16'h276F, 16'h0001,
16'h2770, 16'h0001,
16'h2771, 16'h0001,
16'h2772, 16'h0001,
16'h2773, 16'h0001,
16'h2774, 16'h0001,
16'h2775, 16'h0001,
16'h2776, 16'h0001,
16'h2777, 16'h0001,
16'h2778, 16'h0001,
16'h2779, 16'h0001,
16'h277A, 16'h0001,
16'h277B, 16'h0001,
16'h277C, 16'h0001,
16'h277D, 16'h0001,
16'h277E, 16'h0001,
16'h277F, 16'h0001,
16'h2780, 16'h0001,
16'h2781, 16'h0001,
16'h2782, 16'h0001,
16'h2783, 16'h0001,
16'h2784, 16'h0001,
16'h2785, 16'h0001,
16'h2786, 16'h0001,
16'h2787, 16'h0001,
16'h2788, 16'h0001,
16'h2789, 16'h0001,
16'h278A, 16'h0001,
16'h278B, 16'h0001,
16'h278C, 16'h0001,
16'h278D, 16'h0001,
16'h278E, 16'h0001,
16'h278F, 16'h0001,
16'h2790, 16'h0001,
16'h2791, 16'h0001,
16'h2792, 16'h0001,
16'h2793, 16'h0001,
16'h2794, 16'h0001,
16'h2795, 16'h0001,
16'h2796, 16'h0001,
16'h2797, 16'h0001,
16'h2798, 16'h0001,
16'h2799, 16'h0001,
16'h279A, 16'h0001,
16'h279B, 16'h0001,
16'h279C, 16'h0001,
16'h279D, 16'h0001,
16'h279E, 16'h0001,
16'h279F, 16'h0001,
16'h27A0, 16'h0001,
16'h27A1, 16'h0001,
16'h27A2, 16'h0001,
16'h27A3, 16'h0001,
16'h27A4, 16'h0001,
16'h27A5, 16'h0001,
16'h27A6, 16'h0001,
16'h27A7, 16'h0001,
16'h27A8, 16'h0001,
16'h27A9, 16'h0001,
16'h27AA, 16'h0001,
16'h27AB, 16'h0001,
16'h27AC, 16'h0001,
16'h27AD, 16'h0001,
16'h27AE, 16'h0001,
16'h27AF, 16'h0001,
16'h27B0, 16'h0001,
16'h27B1, 16'h0001,
16'h27B2, 16'h0001,
16'h27B3, 16'h0001,
16'h27B4, 16'h0001,
16'h27B5, 16'h0001,
16'h27B6, 16'h0001,
16'h27B7, 16'h0001,
16'h27B8, 16'h0001,
16'h27B9, 16'h0001,
16'h27BA, 16'h0001,
16'h27BB, 16'h0001,
16'h27BC, 16'h0001,
16'h27BD, 16'h0001,
16'h27BE, 16'h0001,
16'h27BF, 16'h0001,
16'h27C0, 16'h0055,
16'h27C1, 16'h0055,
16'h27C2, 16'h0055,
16'h27C3, 16'h0055,
16'h27C4, 16'h0055,
16'h27C5, 16'h0055,
16'h27C6, 16'h0055,
16'h27C7, 16'h0055,
16'h27C8, 16'h0055,
16'h27C9, 16'h0055,
16'h27CA, 16'h0055,
16'h27CB, 16'h0055,
16'h27CC, 16'h0055,
16'h27CD, 16'h0055,
16'h27CE, 16'h0055,
16'h27CF, 16'h0055,
16'h27D0, 16'h0055,
16'h27D1, 16'h0055,
16'h27D2, 16'h0055,
16'h27D3, 16'h0055,
16'h27D4, 16'h0055,
16'h27D5, 16'h0055,
16'h27D6, 16'h0055,
16'h27D7, 16'h0055,
16'h27D8, 16'h0055,
16'h27D9, 16'h0055,
16'h27DA, 16'h0055,
16'h27DB, 16'h0055,
16'h27DC, 16'h0055,
16'h27DD, 16'h0055,
16'h27DE, 16'h0055,
16'h27DF, 16'h0055,
16'h27E0, 16'h0055,
16'h27E1, 16'h0055,
16'h27E2, 16'h0055,
16'h27E3, 16'h0055,
16'h27E4, 16'h0055,
16'h27E5, 16'h0055,
16'h27E6, 16'h0055,
16'h27E7, 16'h0055,
16'h27E8, 16'h0055,
16'h27E9, 16'h0055,
16'h27EA, 16'h0055,
16'h27EB, 16'h0055,
16'h27EC, 16'h0055,
16'h27ED, 16'h0055,
16'h27EE, 16'h0055,
16'h27EF, 16'h0055,
16'h27F0, 16'h0055,
16'h27F1, 16'h0055,
16'h27F2, 16'h0055,
16'h27F3, 16'h0055,
16'h27F4, 16'h0055,
16'h27F5, 16'h0055,
16'h27F6, 16'h0055,
16'h27F7, 16'h0055,
16'h27F8, 16'h0055,
16'h27F9, 16'h0055,
16'h27FA, 16'h0055,
16'h27FB, 16'h0055,
16'h27FC, 16'h0055,
16'h27FD, 16'h0055,
16'h27FE, 16'h0055,
16'h27FF, 16'h0055,
16'h2800, 16'h0002,
16'h2801, 16'h0002,
16'h2802, 16'h0002,
16'h2803, 16'h0002,
16'h2804, 16'h0002,
16'h2805, 16'h0002,
16'h2806, 16'h0002,
16'h2807, 16'h0002,
16'h2808, 16'h0002,
16'h2809, 16'h0002,
16'h280A, 16'h0002,
16'h280B, 16'h0002,
16'h280C, 16'h0002,
16'h280D, 16'h0002,
16'h280E, 16'h0002,
16'h280F, 16'h0002,
16'h2810, 16'h0002,
16'h2811, 16'h0002,
16'h2812, 16'h0002,
16'h2813, 16'h0002,
16'h2814, 16'h0002,
16'h2815, 16'h0002,
16'h2816, 16'h0002,
16'h2817, 16'h0002,
16'h2818, 16'h0002,
16'h2819, 16'h0002,
16'h281A, 16'h0002,
16'h281B, 16'h0002,
16'h281C, 16'h0002,
16'h281D, 16'h0002,
16'h281E, 16'h0002,
16'h281F, 16'h0002,
16'h2820, 16'h0002,
16'h2821, 16'h0002,
16'h2822, 16'h0002,
16'h2823, 16'h0002,
16'h2824, 16'h0002,
16'h2825, 16'h0002,
16'h2826, 16'h0002,
16'h2827, 16'h0002,
16'h2828, 16'h0002,
16'h2829, 16'h0002,
16'h282A, 16'h0002,
16'h282B, 16'h0002,
16'h282C, 16'h0002,
16'h282D, 16'h0002,
16'h282E, 16'h0002,
16'h282F, 16'h0002,
16'h2830, 16'h0002,
16'h2831, 16'h0002,
16'h2832, 16'h0002,
16'h2833, 16'h0002,
16'h2834, 16'h0002,
16'h2835, 16'h0002,
16'h2836, 16'h0002,
16'h2837, 16'h0002,
16'h2838, 16'h0002,
16'h2839, 16'h0002,
16'h283A, 16'h0002,
16'h283B, 16'h0002,
16'h283C, 16'h0002,
16'h283D, 16'h0002,
16'h283E, 16'h0002,
16'h283F, 16'h0002,
16'h2840, 16'h0002,
16'h2841, 16'h0002,
16'h2842, 16'h0002,
16'h2843, 16'h0002,
16'h2844, 16'h0002,
16'h2845, 16'h0002,
16'h2846, 16'h0002,
16'h2847, 16'h0002,
16'h2848, 16'h0002,
16'h2849, 16'h0002,
16'h284A, 16'h0002,
16'h284B, 16'h0002,
16'h284C, 16'h0002,
16'h284D, 16'h0002,
16'h284E, 16'h0002,
16'h284F, 16'h0002,
16'h2850, 16'h0002,
16'h2851, 16'h0002,
16'h2852, 16'h0002,
16'h2853, 16'h0002,
16'h2854, 16'h0002,
16'h2855, 16'h0002,
16'h2856, 16'h0002,
16'h2857, 16'h0002,
16'h2858, 16'h0002,
16'h2859, 16'h0002,
16'h285A, 16'h0002,
16'h285B, 16'h0002,
16'h285C, 16'h0002,
16'h285D, 16'h0002,
16'h285E, 16'h0002,
16'h285F, 16'h0002,
16'h2860, 16'h0002,
16'h2861, 16'h0002,
16'h2862, 16'h0002,
16'h2863, 16'h0002,
16'h2864, 16'h0002,
16'h2865, 16'h0002,
16'h2866, 16'h0002,
16'h2867, 16'h0002,
16'h2868, 16'h0002,
16'h2869, 16'h0002,
16'h286A, 16'h0002,
16'h286B, 16'h0002,
16'h286C, 16'h0002,
16'h286D, 16'h0002,
16'h286E, 16'h0002,
16'h286F, 16'h0002,
16'h2870, 16'h0002,
16'h2871, 16'h0002,
16'h2872, 16'h0002,
16'h2873, 16'h0002,
16'h2874, 16'h0002,
16'h2875, 16'h0002,
16'h2876, 16'h0002,
16'h2877, 16'h0002,
16'h2878, 16'h0002,
16'h2879, 16'h0002,
16'h287A, 16'h0002,
16'h287B, 16'h0002,
16'h287C, 16'h0002,
16'h287D, 16'h0002,
16'h287E, 16'h0002,
16'h287F, 16'h0002,
16'h2880, 16'h0002,
16'h2881, 16'h0002,
16'h2882, 16'h0002,
16'h2883, 16'h0002,
16'h2884, 16'h0002,
16'h2885, 16'h0002,
16'h2886, 16'h0002,
16'h2887, 16'h0002,
16'h2888, 16'h0002,
16'h2889, 16'h0002,
16'h288A, 16'h0002,
16'h288B, 16'h0002,
16'h288C, 16'h0002,
16'h288D, 16'h0002,
16'h288E, 16'h0002,
16'h288F, 16'h0002,
16'h2890, 16'h0002,
16'h2891, 16'h0002,
16'h2892, 16'h0002,
16'h2893, 16'h0002,
16'h2894, 16'h0002,
16'h2895, 16'h0002,
16'h2896, 16'h0002,
16'h2897, 16'h0002,
16'h2898, 16'h0002,
16'h2899, 16'h0002,
16'h289A, 16'h0002,
16'h289B, 16'h0002,
16'h289C, 16'h0002,
16'h289D, 16'h0002,
16'h289E, 16'h0002,
16'h289F, 16'h0002,
16'h28A0, 16'h0002,
16'h28A1, 16'h0002,
16'h28A2, 16'h0002,
16'h28A3, 16'h0002,
16'h28A4, 16'h0002,
16'h28A5, 16'h0002,
16'h28A6, 16'h0002,
16'h28A7, 16'h0002,
16'h28A8, 16'h0002,
16'h28A9, 16'h0002,
16'h28AA, 16'h0002,
16'h28AB, 16'h0002,
16'h28AC, 16'h0002,
16'h28AD, 16'h0002,
16'h28AE, 16'h0002,
16'h28AF, 16'h0002,
16'h28B0, 16'h0002,
16'h28B1, 16'h0002,
16'h28B2, 16'h0002,
16'h28B3, 16'h0002,
16'h28B4, 16'h0002,
16'h28B5, 16'h0002,
16'h28B6, 16'h0002,
16'h28B7, 16'h0002,
16'h28B8, 16'h0002,
16'h28B9, 16'h0002,
16'h28BA, 16'h0002,
16'h28BB, 16'h0002,
16'h28BC, 16'h0002,
16'h28BD, 16'h0002,
16'h28BE, 16'h0002,
16'h28BF, 16'h0002,
16'h28C0, 16'h0002,
16'h28C1, 16'h0002,
16'h28C2, 16'h0002,
16'h28C3, 16'h0002,
16'h28C4, 16'h0002,
16'h28C5, 16'h0002,
16'h28C6, 16'h0002,
16'h28C7, 16'h0002,
16'h28C8, 16'h0002,
16'h28C9, 16'h0002,
16'h28CA, 16'h0002,
16'h28CB, 16'h0002,
16'h28CC, 16'h0002,
16'h28CD, 16'h0002,
16'h28CE, 16'h0002,
16'h28CF, 16'h0002,
16'h28D0, 16'h0002,
16'h28D1, 16'h0002,
16'h28D2, 16'h0002,
16'h28D3, 16'h0002,
16'h28D4, 16'h0002,
16'h28D5, 16'h0002,
16'h28D6, 16'h0002,
16'h28D7, 16'h0002,
16'h28D8, 16'h0002,
16'h28D9, 16'h0002,
16'h28DA, 16'h0002,
16'h28DB, 16'h0002,
16'h28DC, 16'h0002,
16'h28DD, 16'h0002,
16'h28DE, 16'h0002,
16'h28DF, 16'h0002,
16'h28E0, 16'h0002,
16'h28E1, 16'h0002,
16'h28E2, 16'h0002,
16'h28E3, 16'h0002,
16'h28E4, 16'h0002,
16'h28E5, 16'h0002,
16'h28E6, 16'h0002,
16'h28E7, 16'h0002,
16'h28E8, 16'h0002,
16'h28E9, 16'h0002,
16'h28EA, 16'h0002,
16'h28EB, 16'h0002,
16'h28EC, 16'h0002,
16'h28ED, 16'h0002,
16'h28EE, 16'h0002,
16'h28EF, 16'h0002,
16'h28F0, 16'h0002,
16'h28F1, 16'h0002,
16'h28F2, 16'h0002,
16'h28F3, 16'h0002,
16'h28F4, 16'h0002,
16'h28F5, 16'h0002,
16'h28F6, 16'h0002,
16'h28F7, 16'h0002,
16'h28F8, 16'h0002,
16'h28F9, 16'h0002,
16'h28FA, 16'h0002,
16'h28FB, 16'h0002,
16'h28FC, 16'h0002,
16'h28FD, 16'h0002,
16'h28FE, 16'h0002,
16'h28FF, 16'h0002,
16'h2900, 16'h0002,
16'h2901, 16'h0002,
16'h2902, 16'h0002,
16'h2903, 16'h0002,
16'h2904, 16'h0002,
16'h2905, 16'h0002,
16'h2906, 16'h0002,
16'h2907, 16'h0002,
16'h2908, 16'h0002,
16'h2909, 16'h0002,
16'h290A, 16'h0002,
16'h290B, 16'h0002,
16'h290C, 16'h0002,
16'h290D, 16'h0002,
16'h290E, 16'h0002,
16'h290F, 16'h0002,
16'h2910, 16'h0002,
16'h2911, 16'h0002,
16'h2912, 16'h0002,
16'h2913, 16'h0002,
16'h2914, 16'h0002,
16'h2915, 16'h0002,
16'h2916, 16'h0002,
16'h2917, 16'h0002,
16'h2918, 16'h0002,
16'h2919, 16'h0002,
16'h291A, 16'h0002,
16'h291B, 16'h0002,
16'h291C, 16'h0002,
16'h291D, 16'h0002,
16'h291E, 16'h0002,
16'h291F, 16'h0002,
16'h2920, 16'h0002,
16'h2921, 16'h0002,
16'h2922, 16'h0002,
16'h2923, 16'h0002,
16'h2924, 16'h0002,
16'h2925, 16'h0002,
16'h2926, 16'h0002,
16'h2927, 16'h0002,
16'h2928, 16'h0002,
16'h2929, 16'h0002,
16'h292A, 16'h0002,
16'h292B, 16'h0002,
16'h292C, 16'h0002,
16'h292D, 16'h0002,
16'h292E, 16'h0002,
16'h292F, 16'h0002,
16'h2930, 16'h0002,
16'h2931, 16'h0002,
16'h2932, 16'h0002,
16'h2933, 16'h0002,
16'h2934, 16'h0002,
16'h2935, 16'h0002,
16'h2936, 16'h0002,
16'h2937, 16'h0002,
16'h2938, 16'h0002,
16'h2939, 16'h0002,
16'h293A, 16'h0002,
16'h293B, 16'h0002,
16'h293C, 16'h0002,
16'h293D, 16'h0002,
16'h293E, 16'h0002,
16'h293F, 16'h0002,
16'h2940, 16'h0002,
16'h2941, 16'h0002,
16'h2942, 16'h0002,
16'h2943, 16'h0002,
16'h2944, 16'h0002,
16'h2945, 16'h0002,
16'h2946, 16'h0002,
16'h2947, 16'h0002,
16'h2948, 16'h0002,
16'h2949, 16'h0002,
16'h294A, 16'h0002,
16'h294B, 16'h0002,
16'h294C, 16'h0002,
16'h294D, 16'h0002,
16'h294E, 16'h0002,
16'h294F, 16'h0002,
16'h2950, 16'h0002,
16'h2951, 16'h0002,
16'h2952, 16'h0002,
16'h2953, 16'h0002,
16'h2954, 16'h0002,
16'h2955, 16'h0002,
16'h2956, 16'h0002,
16'h2957, 16'h0002,
16'h2958, 16'h0002,
16'h2959, 16'h0002,
16'h295A, 16'h0002,
16'h295B, 16'h0002,
16'h295C, 16'h0002,
16'h295D, 16'h0002,
16'h295E, 16'h0002,
16'h295F, 16'h0002,
16'h2960, 16'h0002,
16'h2961, 16'h0002,
16'h2962, 16'h0002,
16'h2963, 16'h0002,
16'h2964, 16'h0002,
16'h2965, 16'h0002,
16'h2966, 16'h0002,
16'h2967, 16'h0002,
16'h2968, 16'h0002,
16'h2969, 16'h0002,
16'h296A, 16'h0002,
16'h296B, 16'h0002,
16'h296C, 16'h0002,
16'h296D, 16'h0002,
16'h296E, 16'h0002,
16'h296F, 16'h0002,
16'h2970, 16'h0002,
16'h2971, 16'h0002,
16'h2972, 16'h0002,
16'h2973, 16'h0002,
16'h2974, 16'h0002,
16'h2975, 16'h0002,
16'h2976, 16'h0002,
16'h2977, 16'h0002,
16'h2978, 16'h0002,
16'h2979, 16'h0002,
16'h297A, 16'h0002,
16'h297B, 16'h0002,
16'h297C, 16'h0002,
16'h297D, 16'h0002,
16'h297E, 16'h0002,
16'h297F, 16'h0002,
16'h2980, 16'h0002,
16'h2981, 16'h0002,
16'h2982, 16'h0002,
16'h2983, 16'h0002,
16'h2984, 16'h0002,
16'h2985, 16'h0002,
16'h2986, 16'h0002,
16'h2987, 16'h0002,
16'h2988, 16'h0002,
16'h2989, 16'h0002,
16'h298A, 16'h0002,
16'h298B, 16'h0002,
16'h298C, 16'h0002,
16'h298D, 16'h0002,
16'h298E, 16'h0002,
16'h298F, 16'h0002,
16'h2990, 16'h0002,
16'h2991, 16'h0002,
16'h2992, 16'h0002,
16'h2993, 16'h0002,
16'h2994, 16'h0002,
16'h2995, 16'h0002,
16'h2996, 16'h0002,
16'h2997, 16'h0002,
16'h2998, 16'h0002,
16'h2999, 16'h0002,
16'h299A, 16'h0002,
16'h299B, 16'h0002,
16'h299C, 16'h0002,
16'h299D, 16'h0002,
16'h299E, 16'h0002,
16'h299F, 16'h0002,
16'h29A0, 16'h0002,
16'h29A1, 16'h0002,
16'h29A2, 16'h0002,
16'h29A3, 16'h0002,
16'h29A4, 16'h0002,
16'h29A5, 16'h0002,
16'h29A6, 16'h0002,
16'h29A7, 16'h0002,
16'h29A8, 16'h0002,
16'h29A9, 16'h0002,
16'h29AA, 16'h0002,
16'h29AB, 16'h0002,
16'h29AC, 16'h0002,
16'h29AD, 16'h0002,
16'h29AE, 16'h0002,
16'h29AF, 16'h0002,
16'h29B0, 16'h0002,
16'h29B1, 16'h0002,
16'h29B2, 16'h0002,
16'h29B3, 16'h0002,
16'h29B4, 16'h0002,
16'h29B5, 16'h0002,
16'h29B6, 16'h0002,
16'h29B7, 16'h0002,
16'h29B8, 16'h0002,
16'h29B9, 16'h0002,
16'h29BA, 16'h0002,
16'h29BB, 16'h0002,
16'h29BC, 16'h0002,
16'h29BD, 16'h0002,
16'h29BE, 16'h0002,
16'h29BF, 16'h0002,
16'h29C0, 16'h0002,
16'h29C1, 16'h0002,
16'h29C2, 16'h0002,
16'h29C3, 16'h0002,
16'h29C4, 16'h0002,
16'h29C5, 16'h0002,
16'h29C6, 16'h0002,
16'h29C7, 16'h0002,
16'h29C8, 16'h0002,
16'h29C9, 16'h0002,
16'h29CA, 16'h0002,
16'h29CB, 16'h0002,
16'h29CC, 16'h0002,
16'h29CD, 16'h0002,
16'h29CE, 16'h0002,
16'h29CF, 16'h0002,
16'h29D0, 16'h0002,
16'h29D1, 16'h0002,
16'h29D2, 16'h0002,
16'h29D3, 16'h0002,
16'h29D4, 16'h0002,
16'h29D5, 16'h0002,
16'h29D6, 16'h0002,
16'h29D7, 16'h0002,
16'h29D8, 16'h0002,
16'h29D9, 16'h0002,
16'h29DA, 16'h0002,
16'h29DB, 16'h0002,
16'h29DC, 16'h0002,
16'h29DD, 16'h0002,
16'h29DE, 16'h0002,
16'h29DF, 16'h0002,
16'h29E0, 16'h0002,
16'h29E1, 16'h0002,
16'h29E2, 16'h0002,
16'h29E3, 16'h0002,
16'h29E4, 16'h0002,
16'h29E5, 16'h0002,
16'h29E6, 16'h0002,
16'h29E7, 16'h0002,
16'h29E8, 16'h0002,
16'h29E9, 16'h0002,
16'h29EA, 16'h0002,
16'h29EB, 16'h0002,
16'h29EC, 16'h0002,
16'h29ED, 16'h0002,
16'h29EE, 16'h0002,
16'h29EF, 16'h0002,
16'h29F0, 16'h0002,
16'h29F1, 16'h0002,
16'h29F2, 16'h0002,
16'h29F3, 16'h0002,
16'h29F4, 16'h0002,
16'h29F5, 16'h0002,
16'h29F6, 16'h0002,
16'h29F7, 16'h0002,
16'h29F8, 16'h0002,
16'h29F9, 16'h0002,
16'h29FA, 16'h0002,
16'h29FB, 16'h0002,
16'h29FC, 16'h0002,
16'h29FD, 16'h0002,
16'h29FE, 16'h0002,
16'h29FF, 16'h0002,
16'h2A00, 16'h0002,
16'h2A01, 16'h0002,
16'h2A02, 16'h0002,
16'h2A03, 16'h0002,
16'h2A04, 16'h0002,
16'h2A05, 16'h0002,
16'h2A06, 16'h0002,
16'h2A07, 16'h0002,
16'h2A08, 16'h0002,
16'h2A09, 16'h0002,
16'h2A0A, 16'h0002,
16'h2A0B, 16'h0002,
16'h2A0C, 16'h0002,
16'h2A0D, 16'h0002,
16'h2A0E, 16'h0002,
16'h2A0F, 16'h0002,
16'h2A10, 16'h0002,
16'h2A11, 16'h0002,
16'h2A12, 16'h0002,
16'h2A13, 16'h0002,
16'h2A14, 16'h0002,
16'h2A15, 16'h0002,
16'h2A16, 16'h0002,
16'h2A17, 16'h0002,
16'h2A18, 16'h0002,
16'h2A19, 16'h0002,
16'h2A1A, 16'h0002,
16'h2A1B, 16'h0002,
16'h2A1C, 16'h0002,
16'h2A1D, 16'h0002,
16'h2A1E, 16'h0002,
16'h2A1F, 16'h0002,
16'h2A20, 16'h0002,
16'h2A21, 16'h0002,
16'h2A22, 16'h0002,
16'h2A23, 16'h0002,
16'h2A24, 16'h0002,
16'h2A25, 16'h0002,
16'h2A26, 16'h0002,
16'h2A27, 16'h0002,
16'h2A28, 16'h0002,
16'h2A29, 16'h0002,
16'h2A2A, 16'h0002,
16'h2A2B, 16'h0002,
16'h2A2C, 16'h0002,
16'h2A2D, 16'h0002,
16'h2A2E, 16'h0002,
16'h2A2F, 16'h0002,
16'h2A30, 16'h0002,
16'h2A31, 16'h0002,
16'h2A32, 16'h0002,
16'h2A33, 16'h0002,
16'h2A34, 16'h0002,
16'h2A35, 16'h0002,
16'h2A36, 16'h0002,
16'h2A37, 16'h0002,
16'h2A38, 16'h0002,
16'h2A39, 16'h0002,
16'h2A3A, 16'h0002,
16'h2A3B, 16'h0002,
16'h2A3C, 16'h0002,
16'h2A3D, 16'h0002,
16'h2A3E, 16'h0002,
16'h2A3F, 16'h0002,
16'h2A40, 16'h0002,
16'h2A41, 16'h0002,
16'h2A42, 16'h0002,
16'h2A43, 16'h0002,
16'h2A44, 16'h0002,
16'h2A45, 16'h0002,
16'h2A46, 16'h0002,
16'h2A47, 16'h0002,
16'h2A48, 16'h0002,
16'h2A49, 16'h0002,
16'h2A4A, 16'h0002,
16'h2A4B, 16'h0002,
16'h2A4C, 16'h0002,
16'h2A4D, 16'h0002,
16'h2A4E, 16'h0002,
16'h2A4F, 16'h0002,
16'h2A50, 16'h0002,
16'h2A51, 16'h0002,
16'h2A52, 16'h0002,
16'h2A53, 16'h0002,
16'h2A54, 16'h0002,
16'h2A55, 16'h0002,
16'h2A56, 16'h0002,
16'h2A57, 16'h0002,
16'h2A58, 16'h0002,
16'h2A59, 16'h0002,
16'h2A5A, 16'h0002,
16'h2A5B, 16'h0002,
16'h2A5C, 16'h0002,
16'h2A5D, 16'h0002,
16'h2A5E, 16'h0002,
16'h2A5F, 16'h0002,
16'h2A60, 16'h0002,
16'h2A61, 16'h0002,
16'h2A62, 16'h0002,
16'h2A63, 16'h0002,
16'h2A64, 16'h0002,
16'h2A65, 16'h0002,
16'h2A66, 16'h0002,
16'h2A67, 16'h0002,
16'h2A68, 16'h0002,
16'h2A69, 16'h0002,
16'h2A6A, 16'h0002,
16'h2A6B, 16'h0002,
16'h2A6C, 16'h0002,
16'h2A6D, 16'h0002,
16'h2A6E, 16'h0002,
16'h2A6F, 16'h0002,
16'h2A70, 16'h0002,
16'h2A71, 16'h0002,
16'h2A72, 16'h0002,
16'h2A73, 16'h0002,
16'h2A74, 16'h0002,
16'h2A75, 16'h0002,
16'h2A76, 16'h0002,
16'h2A77, 16'h0002,
16'h2A78, 16'h0002,
16'h2A79, 16'h0002,
16'h2A7A, 16'h0002,
16'h2A7B, 16'h0002,
16'h2A7C, 16'h0002,
16'h2A7D, 16'h0002,
16'h2A7E, 16'h0002,
16'h2A7F, 16'h0002,
16'h2A80, 16'h0002,
16'h2A81, 16'h0002,
16'h2A82, 16'h0002,
16'h2A83, 16'h0002,
16'h2A84, 16'h0002,
16'h2A85, 16'h0002,
16'h2A86, 16'h0002,
16'h2A87, 16'h0002,
16'h2A88, 16'h0002,
16'h2A89, 16'h0002,
16'h2A8A, 16'h0002,
16'h2A8B, 16'h0002,
16'h2A8C, 16'h0002,
16'h2A8D, 16'h0002,
16'h2A8E, 16'h0002,
16'h2A8F, 16'h0002,
16'h2A90, 16'h0002,
16'h2A91, 16'h0002,
16'h2A92, 16'h0002,
16'h2A93, 16'h0002,
16'h2A94, 16'h0002,
16'h2A95, 16'h0002,
16'h2A96, 16'h0002,
16'h2A97, 16'h0002,
16'h2A98, 16'h0002,
16'h2A99, 16'h0002,
16'h2A9A, 16'h0002,
16'h2A9B, 16'h0002,
16'h2A9C, 16'h0002,
16'h2A9D, 16'h0002,
16'h2A9E, 16'h0002,
16'h2A9F, 16'h0002,
16'h2AA0, 16'h0002,
16'h2AA1, 16'h0002,
16'h2AA2, 16'h0002,
16'h2AA3, 16'h0002,
16'h2AA4, 16'h0002,
16'h2AA5, 16'h0002,
16'h2AA6, 16'h0002,
16'h2AA7, 16'h0002,
16'h2AA8, 16'h0002,
16'h2AA9, 16'h0002,
16'h2AAA, 16'h0002,
16'h2AAB, 16'h0002,
16'h2AAC, 16'h0002,
16'h2AAD, 16'h0002,
16'h2AAE, 16'h0002,
16'h2AAF, 16'h0002,
16'h2AB0, 16'h0002,
16'h2AB1, 16'h0002,
16'h2AB2, 16'h0002,
16'h2AB3, 16'h0002,
16'h2AB4, 16'h0002,
16'h2AB5, 16'h0002,
16'h2AB6, 16'h0002,
16'h2AB7, 16'h0002,
16'h2AB8, 16'h0002,
16'h2AB9, 16'h0002,
16'h2ABA, 16'h0002,
16'h2ABB, 16'h0002,
16'h2ABC, 16'h0002,
16'h2ABD, 16'h0002,
16'h2ABE, 16'h0002,
16'h2ABF, 16'h0002,
16'h2AC0, 16'h0002,
16'h2AC1, 16'h0002,
16'h2AC2, 16'h0002,
16'h2AC3, 16'h0002,
16'h2AC4, 16'h0002,
16'h2AC5, 16'h0002,
16'h2AC6, 16'h0002,
16'h2AC7, 16'h0002,
16'h2AC8, 16'h0002,
16'h2AC9, 16'h0002,
16'h2ACA, 16'h0002,
16'h2ACB, 16'h0002,
16'h2ACC, 16'h0002,
16'h2ACD, 16'h0002,
16'h2ACE, 16'h0002,
16'h2ACF, 16'h0002,
16'h2AD0, 16'h0002,
16'h2AD1, 16'h0002,
16'h2AD2, 16'h0002,
16'h2AD3, 16'h0002,
16'h2AD4, 16'h0002,
16'h2AD5, 16'h0002,
16'h2AD6, 16'h0002,
16'h2AD7, 16'h0002,
16'h2AD8, 16'h0002,
16'h2AD9, 16'h0002,
16'h2ADA, 16'h0002,
16'h2ADB, 16'h0002,
16'h2ADC, 16'h0002,
16'h2ADD, 16'h0002,
16'h2ADE, 16'h0002,
16'h2ADF, 16'h0002,
16'h2AE0, 16'h0002,
16'h2AE1, 16'h0002,
16'h2AE2, 16'h0002,
16'h2AE3, 16'h0002,
16'h2AE4, 16'h0002,
16'h2AE5, 16'h0002,
16'h2AE6, 16'h0002,
16'h2AE7, 16'h0002,
16'h2AE8, 16'h0002,
16'h2AE9, 16'h0002,
16'h2AEA, 16'h0002,
16'h2AEB, 16'h0002,
16'h2AEC, 16'h0002,
16'h2AED, 16'h0002,
16'h2AEE, 16'h0002,
16'h2AEF, 16'h0002,
16'h2AF0, 16'h0002,
16'h2AF1, 16'h0002,
16'h2AF2, 16'h0002,
16'h2AF3, 16'h0002,
16'h2AF4, 16'h0002,
16'h2AF5, 16'h0002,
16'h2AF6, 16'h0002,
16'h2AF7, 16'h0002,
16'h2AF8, 16'h0002,
16'h2AF9, 16'h0002,
16'h2AFA, 16'h0002,
16'h2AFB, 16'h0002,
16'h2AFC, 16'h0002,
16'h2AFD, 16'h0002,
16'h2AFE, 16'h0002,
16'h2AFF, 16'h0002,
16'h2B00, 16'h0002,
16'h2B01, 16'h0002,
16'h2B02, 16'h0002,
16'h2B03, 16'h0002,
16'h2B04, 16'h0002,
16'h2B05, 16'h0002,
16'h2B06, 16'h0002,
16'h2B07, 16'h0002,
16'h2B08, 16'h0002,
16'h2B09, 16'h0002,
16'h2B0A, 16'h0002,
16'h2B0B, 16'h0002,
16'h2B0C, 16'h0002,
16'h2B0D, 16'h0002,
16'h2B0E, 16'h0002,
16'h2B0F, 16'h0002,
16'h2B10, 16'h0002,
16'h2B11, 16'h0002,
16'h2B12, 16'h0002,
16'h2B13, 16'h0002,
16'h2B14, 16'h0002,
16'h2B15, 16'h0002,
16'h2B16, 16'h0002,
16'h2B17, 16'h0002,
16'h2B18, 16'h0002,
16'h2B19, 16'h0002,
16'h2B1A, 16'h0002,
16'h2B1B, 16'h0002,
16'h2B1C, 16'h0002,
16'h2B1D, 16'h0002,
16'h2B1E, 16'h0002,
16'h2B1F, 16'h0002,
16'h2B20, 16'h0002,
16'h2B21, 16'h0002,
16'h2B22, 16'h0002,
16'h2B23, 16'h0002,
16'h2B24, 16'h0002,
16'h2B25, 16'h0002,
16'h2B26, 16'h0002,
16'h2B27, 16'h0002,
16'h2B28, 16'h0002,
16'h2B29, 16'h0002,
16'h2B2A, 16'h0002,
16'h2B2B, 16'h0002,
16'h2B2C, 16'h0002,
16'h2B2D, 16'h0002,
16'h2B2E, 16'h0002,
16'h2B2F, 16'h0002,
16'h2B30, 16'h0002,
16'h2B31, 16'h0002,
16'h2B32, 16'h0002,
16'h2B33, 16'h0002,
16'h2B34, 16'h0002,
16'h2B35, 16'h0002,
16'h2B36, 16'h0002,
16'h2B37, 16'h0002,
16'h2B38, 16'h0002,
16'h2B39, 16'h0002,
16'h2B3A, 16'h0002,
16'h2B3B, 16'h0002,
16'h2B3C, 16'h0002,
16'h2B3D, 16'h0002,
16'h2B3E, 16'h0002,
16'h2B3F, 16'h0002,
16'h2B40, 16'h0002,
16'h2B41, 16'h0002,
16'h2B42, 16'h0002,
16'h2B43, 16'h0002,
16'h2B44, 16'h0002,
16'h2B45, 16'h0002,
16'h2B46, 16'h0002,
16'h2B47, 16'h0002,
16'h2B48, 16'h0002,
16'h2B49, 16'h0002,
16'h2B4A, 16'h0002,
16'h2B4B, 16'h0002,
16'h2B4C, 16'h0002,
16'h2B4D, 16'h0002,
16'h2B4E, 16'h0002,
16'h2B4F, 16'h0002,
16'h2B50, 16'h0002,
16'h2B51, 16'h0002,
16'h2B52, 16'h0002,
16'h2B53, 16'h0002,
16'h2B54, 16'h0002,
16'h2B55, 16'h0002,
16'h2B56, 16'h0002,
16'h2B57, 16'h0002,
16'h2B58, 16'h0002,
16'h2B59, 16'h0002,
16'h2B5A, 16'h0002,
16'h2B5B, 16'h0002,
16'h2B5C, 16'h0002,
16'h2B5D, 16'h0002,
16'h2B5E, 16'h0002,
16'h2B5F, 16'h0002,
16'h2B60, 16'h0002,
16'h2B61, 16'h0002,
16'h2B62, 16'h0002,
16'h2B63, 16'h0002,
16'h2B64, 16'h0002,
16'h2B65, 16'h0002,
16'h2B66, 16'h0002,
16'h2B67, 16'h0002,
16'h2B68, 16'h0002,
16'h2B69, 16'h0002,
16'h2B6A, 16'h0002,
16'h2B6B, 16'h0002,
16'h2B6C, 16'h0002,
16'h2B6D, 16'h0002,
16'h2B6E, 16'h0002,
16'h2B6F, 16'h0002,
16'h2B70, 16'h0002,
16'h2B71, 16'h0002,
16'h2B72, 16'h0002,
16'h2B73, 16'h0002,
16'h2B74, 16'h0002,
16'h2B75, 16'h0002,
16'h2B76, 16'h0002,
16'h2B77, 16'h0002,
16'h2B78, 16'h0002,
16'h2B79, 16'h0002,
16'h2B7A, 16'h0002,
16'h2B7B, 16'h0002,
16'h2B7C, 16'h0002,
16'h2B7D, 16'h0002,
16'h2B7E, 16'h0002,
16'h2B7F, 16'h0002,
16'h2B80, 16'h0002,
16'h2B81, 16'h0002,
16'h2B82, 16'h0002,
16'h2B83, 16'h0002,
16'h2B84, 16'h0002,
16'h2B85, 16'h0002,
16'h2B86, 16'h0002,
16'h2B87, 16'h0002,
16'h2B88, 16'h0002,
16'h2B89, 16'h0002,
16'h2B8A, 16'h0002,
16'h2B8B, 16'h0002,
16'h2B8C, 16'h0002,
16'h2B8D, 16'h0002,
16'h2B8E, 16'h0002,
16'h2B8F, 16'h0002,
16'h2B90, 16'h0002,
16'h2B91, 16'h0002,
16'h2B92, 16'h0002,
16'h2B93, 16'h0002,
16'h2B94, 16'h0002,
16'h2B95, 16'h0002,
16'h2B96, 16'h0002,
16'h2B97, 16'h0002,
16'h2B98, 16'h0002,
16'h2B99, 16'h0002,
16'h2B9A, 16'h0002,
16'h2B9B, 16'h0002,
16'h2B9C, 16'h0002,
16'h2B9D, 16'h0002,
16'h2B9E, 16'h0002,
16'h2B9F, 16'h0002,
16'h2BA0, 16'h0002,
16'h2BA1, 16'h0002,
16'h2BA2, 16'h0002,
16'h2BA3, 16'h0002,
16'h2BA4, 16'h0002,
16'h2BA5, 16'h0002,
16'h2BA6, 16'h0002,
16'h2BA7, 16'h0002,
16'h2BA8, 16'h0002,
16'h2BA9, 16'h0002,
16'h2BAA, 16'h0002,
16'h2BAB, 16'h0002,
16'h2BAC, 16'h0002,
16'h2BAD, 16'h0002,
16'h2BAE, 16'h0002,
16'h2BAF, 16'h0002,
16'h2BB0, 16'h0002,
16'h2BB1, 16'h0002,
16'h2BB2, 16'h0002,
16'h2BB3, 16'h0002,
16'h2BB4, 16'h0002,
16'h2BB5, 16'h0002,
16'h2BB6, 16'h0002,
16'h2BB7, 16'h0002,
16'h2BB8, 16'h0002,
16'h2BB9, 16'h0002,
16'h2BBA, 16'h0002,
16'h2BBB, 16'h0002,
16'h2BBC, 16'h0002,
16'h2BBD, 16'h0002,
16'h2BBE, 16'h0002,
16'h2BBF, 16'h0002,
16'h2BC0, 16'h00AA,
16'h2BC1, 16'h00AA,
16'h2BC2, 16'h00AA,
16'h2BC3, 16'h00AA,
16'h2BC4, 16'h00AA,
16'h2BC5, 16'h00AA,
16'h2BC6, 16'h00AA,
16'h2BC7, 16'h00AA,
16'h2BC8, 16'h00AA,
16'h2BC9, 16'h00AA,
16'h2BCA, 16'h00AA,
16'h2BCB, 16'h00AA,
16'h2BCC, 16'h00AA,
16'h2BCD, 16'h00AA,
16'h2BCE, 16'h00AA,
16'h2BCF, 16'h00AA,
16'h2BD0, 16'h00AA,
16'h2BD1, 16'h00AA,
16'h2BD2, 16'h00AA,
16'h2BD3, 16'h00AA,
16'h2BD4, 16'h00AA,
16'h2BD5, 16'h00AA,
16'h2BD6, 16'h00AA,
16'h2BD7, 16'h00AA,
16'h2BD8, 16'h00AA,
16'h2BD9, 16'h00AA,
16'h2BDA, 16'h00AA,
16'h2BDB, 16'h00AA,
16'h2BDC, 16'h00AA,
16'h2BDD, 16'h00AA,
16'h2BDE, 16'h00AA,
16'h2BDF, 16'h00AA,
16'h2BE0, 16'h00AA,
16'h2BE1, 16'h00AA,
16'h2BE2, 16'h00AA,
16'h2BE3, 16'h00AA,
16'h2BE4, 16'h00AA,
16'h2BE5, 16'h00AA,
16'h2BE6, 16'h00AA,
16'h2BE7, 16'h00AA,
16'h2BE8, 16'h00AA,
16'h2BE9, 16'h00AA,
16'h2BEA, 16'h00AA,
16'h2BEB, 16'h00AA,
16'h2BEC, 16'h00AA,
16'h2BED, 16'h00AA,
16'h2BEE, 16'h00AA,
16'h2BEF, 16'h00AA,
16'h2BF0, 16'h00AA,
16'h2BF1, 16'h00AA,
16'h2BF2, 16'h00AA,
16'h2BF3, 16'h00AA,
16'h2BF4, 16'h00AA,
16'h2BF5, 16'h00AA,
16'h2BF6, 16'h00AA,
16'h2BF7, 16'h00AA,
16'h2BF8, 16'h00AA,
16'h2BF9, 16'h00AA,
16'h2BFA, 16'h00AA,
16'h2BFB, 16'h00AA,
16'h2BFC, 16'h00AA,
16'h2BFD, 16'h00AA,
16'h2BFE, 16'h00AA,
16'h2BFF, 16'h00AA,
16'h2C00, 16'h0003,
16'h2C01, 16'h0003,
16'h2C02, 16'h0003,
16'h2C03, 16'h0003,
16'h2C04, 16'h0003,
16'h2C05, 16'h0003,
16'h2C06, 16'h0003,
16'h2C07, 16'h0003,
16'h2C08, 16'h0003,
16'h2C09, 16'h0003,
16'h2C0A, 16'h0003,
16'h2C0B, 16'h0003,
16'h2C0C, 16'h0003,
16'h2C0D, 16'h0003,
16'h2C0E, 16'h0003,
16'h2C0F, 16'h0003,
16'h2C10, 16'h0003,
16'h2C11, 16'h0003,
16'h2C12, 16'h0003,
16'h2C13, 16'h0003,
16'h2C14, 16'h0003,
16'h2C15, 16'h0003,
16'h2C16, 16'h0003,
16'h2C17, 16'h0003,
16'h2C18, 16'h0003,
16'h2C19, 16'h0003,
16'h2C1A, 16'h0003,
16'h2C1B, 16'h0003,
16'h2C1C, 16'h0003,
16'h2C1D, 16'h0003,
16'h2C1E, 16'h0003,
16'h2C1F, 16'h0003,
16'h2C20, 16'h0003,
16'h2C21, 16'h0003,
16'h2C22, 16'h0003,
16'h2C23, 16'h0003,
16'h2C24, 16'h0003,
16'h2C25, 16'h0003,
16'h2C26, 16'h0003,
16'h2C27, 16'h0003,
16'h2C28, 16'h0003,
16'h2C29, 16'h0003,
16'h2C2A, 16'h0003,
16'h2C2B, 16'h0003,
16'h2C2C, 16'h0003,
16'h2C2D, 16'h0003,
16'h2C2E, 16'h0003,
16'h2C2F, 16'h0003,
16'h2C30, 16'h0003,
16'h2C31, 16'h0003,
16'h2C32, 16'h0003,
16'h2C33, 16'h0003,
16'h2C34, 16'h0003,
16'h2C35, 16'h0003,
16'h2C36, 16'h0003,
16'h2C37, 16'h0003,
16'h2C38, 16'h0003,
16'h2C39, 16'h0003,
16'h2C3A, 16'h0003,
16'h2C3B, 16'h0003,
16'h2C3C, 16'h0003,
16'h2C3D, 16'h0003,
16'h2C3E, 16'h0003,
16'h2C3F, 16'h0003,
16'h2C40, 16'h0003,
16'h2C41, 16'h0003,
16'h2C42, 16'h0003,
16'h2C43, 16'h0003,
16'h2C44, 16'h0003,
16'h2C45, 16'h0003,
16'h2C46, 16'h0003,
16'h2C47, 16'h0003,
16'h2C48, 16'h0003,
16'h2C49, 16'h0003,
16'h2C4A, 16'h0003,
16'h2C4B, 16'h0003,
16'h2C4C, 16'h0003,
16'h2C4D, 16'h0003,
16'h2C4E, 16'h0003,
16'h2C4F, 16'h0003,
16'h2C50, 16'h0003,
16'h2C51, 16'h0003,
16'h2C52, 16'h0003,
16'h2C53, 16'h0003,
16'h2C54, 16'h0003,
16'h2C55, 16'h0003,
16'h2C56, 16'h0003,
16'h2C57, 16'h0003,
16'h2C58, 16'h0003,
16'h2C59, 16'h0003,
16'h2C5A, 16'h0003,
16'h2C5B, 16'h0003,
16'h2C5C, 16'h0003,
16'h2C5D, 16'h0003,
16'h2C5E, 16'h0003,
16'h2C5F, 16'h0003,
16'h2C60, 16'h0003,
16'h2C61, 16'h0003,
16'h2C62, 16'h0003,
16'h2C63, 16'h0003,
16'h2C64, 16'h0003,
16'h2C65, 16'h0003,
16'h2C66, 16'h0003,
16'h2C67, 16'h0003,
16'h2C68, 16'h0003,
16'h2C69, 16'h0003,
16'h2C6A, 16'h0003,
16'h2C6B, 16'h0003,
16'h2C6C, 16'h0003,
16'h2C6D, 16'h0003,
16'h2C6E, 16'h0003,
16'h2C6F, 16'h0003,
16'h2C70, 16'h0003,
16'h2C71, 16'h0003,
16'h2C72, 16'h0003,
16'h2C73, 16'h0003,
16'h2C74, 16'h0003,
16'h2C75, 16'h0003,
16'h2C76, 16'h0003,
16'h2C77, 16'h0003,
16'h2C78, 16'h0003,
16'h2C79, 16'h0003,
16'h2C7A, 16'h0003,
16'h2C7B, 16'h0003,
16'h2C7C, 16'h0003,
16'h2C7D, 16'h0003,
16'h2C7E, 16'h0003,
16'h2C7F, 16'h0003,
16'h2C80, 16'h0003,
16'h2C81, 16'h0003,
16'h2C82, 16'h0003,
16'h2C83, 16'h0003,
16'h2C84, 16'h0003,
16'h2C85, 16'h0003,
16'h2C86, 16'h0003,
16'h2C87, 16'h0003,
16'h2C88, 16'h0003,
16'h2C89, 16'h0003,
16'h2C8A, 16'h0003,
16'h2C8B, 16'h0003,
16'h2C8C, 16'h0003,
16'h2C8D, 16'h0003,
16'h2C8E, 16'h0003,
16'h2C8F, 16'h0003,
16'h2C90, 16'h0003,
16'h2C91, 16'h0003,
16'h2C92, 16'h0003,
16'h2C93, 16'h0003,
16'h2C94, 16'h0003,
16'h2C95, 16'h0003,
16'h2C96, 16'h0003,
16'h2C97, 16'h0003,
16'h2C98, 16'h0003,
16'h2C99, 16'h0003,
16'h2C9A, 16'h0003,
16'h2C9B, 16'h0003,
16'h2C9C, 16'h0003,
16'h2C9D, 16'h0003,
16'h2C9E, 16'h0003,
16'h2C9F, 16'h0003,
16'h2CA0, 16'h0003,
16'h2CA1, 16'h0003,
16'h2CA2, 16'h0003,
16'h2CA3, 16'h0003,
16'h2CA4, 16'h0003,
16'h2CA5, 16'h0003,
16'h2CA6, 16'h0003,
16'h2CA7, 16'h0003,
16'h2CA8, 16'h0003,
16'h2CA9, 16'h0003,
16'h2CAA, 16'h0003,
16'h2CAB, 16'h0003,
16'h2CAC, 16'h0003,
16'h2CAD, 16'h0003,
16'h2CAE, 16'h0003,
16'h2CAF, 16'h0003,
16'h2CB0, 16'h0003,
16'h2CB1, 16'h0003,
16'h2CB2, 16'h0003,
16'h2CB3, 16'h0003,
16'h2CB4, 16'h0003,
16'h2CB5, 16'h0003,
16'h2CB6, 16'h0003,
16'h2CB7, 16'h0003,
16'h2CB8, 16'h0003,
16'h2CB9, 16'h0003,
16'h2CBA, 16'h0003,
16'h2CBB, 16'h0003,
16'h2CBC, 16'h0003,
16'h2CBD, 16'h0003,
16'h2CBE, 16'h0003,
16'h2CBF, 16'h0003,
16'h2CC0, 16'h0003,
16'h2CC1, 16'h0003,
16'h2CC2, 16'h0003,
16'h2CC3, 16'h0003,
16'h2CC4, 16'h0003,
16'h2CC5, 16'h0003,
16'h2CC6, 16'h0003,
16'h2CC7, 16'h0003,
16'h2CC8, 16'h0003,
16'h2CC9, 16'h0003,
16'h2CCA, 16'h0003,
16'h2CCB, 16'h0003,
16'h2CCC, 16'h0003,
16'h2CCD, 16'h0003,
16'h2CCE, 16'h0003,
16'h2CCF, 16'h0003,
16'h2CD0, 16'h0003,
16'h2CD1, 16'h0003,
16'h2CD2, 16'h0003,
16'h2CD3, 16'h0003,
16'h2CD4, 16'h0003,
16'h2CD5, 16'h0003,
16'h2CD6, 16'h0003,
16'h2CD7, 16'h0003,
16'h2CD8, 16'h0003,
16'h2CD9, 16'h0003,
16'h2CDA, 16'h0003,
16'h2CDB, 16'h0003,
16'h2CDC, 16'h0003,
16'h2CDD, 16'h0003,
16'h2CDE, 16'h0003,
16'h2CDF, 16'h0003,
16'h2CE0, 16'h0003,
16'h2CE1, 16'h0003,
16'h2CE2, 16'h0003,
16'h2CE3, 16'h0003,
16'h2CE4, 16'h0003,
16'h2CE5, 16'h0003,
16'h2CE6, 16'h0003,
16'h2CE7, 16'h0003,
16'h2CE8, 16'h0003,
16'h2CE9, 16'h0003,
16'h2CEA, 16'h0003,
16'h2CEB, 16'h0003,
16'h2CEC, 16'h0003,
16'h2CED, 16'h0003,
16'h2CEE, 16'h0003,
16'h2CEF, 16'h0003,
16'h2CF0, 16'h0003,
16'h2CF1, 16'h0003,
16'h2CF2, 16'h0003,
16'h2CF3, 16'h0003,
16'h2CF4, 16'h0003,
16'h2CF5, 16'h0003,
16'h2CF6, 16'h0003,
16'h2CF7, 16'h0003,
16'h2CF8, 16'h0003,
16'h2CF9, 16'h0003,
16'h2CFA, 16'h0003,
16'h2CFB, 16'h0003,
16'h2CFC, 16'h0003,
16'h2CFD, 16'h0003,
16'h2CFE, 16'h0003,
16'h2CFF, 16'h0003,
16'h2D00, 16'h0003,
16'h2D01, 16'h0003,
16'h2D02, 16'h0003,
16'h2D03, 16'h0003,
16'h2D04, 16'h0003,
16'h2D05, 16'h0003,
16'h2D06, 16'h0003,
16'h2D07, 16'h0003,
16'h2D08, 16'h0003,
16'h2D09, 16'h0003,
16'h2D0A, 16'h0003,
16'h2D0B, 16'h0003,
16'h2D0C, 16'h0003,
16'h2D0D, 16'h0003,
16'h2D0E, 16'h0003,
16'h2D0F, 16'h0003,
16'h2D10, 16'h0003,
16'h2D11, 16'h0003,
16'h2D12, 16'h0003,
16'h2D13, 16'h0003,
16'h2D14, 16'h0003,
16'h2D15, 16'h0003,
16'h2D16, 16'h0003,
16'h2D17, 16'h0003,
16'h2D18, 16'h0003,
16'h2D19, 16'h0003,
16'h2D1A, 16'h0003,
16'h2D1B, 16'h0003,
16'h2D1C, 16'h0003,
16'h2D1D, 16'h0003,
16'h2D1E, 16'h0003,
16'h2D1F, 16'h0003,
16'h2D20, 16'h0003,
16'h2D21, 16'h0003,
16'h2D22, 16'h0003,
16'h2D23, 16'h0003,
16'h2D24, 16'h0003,
16'h2D25, 16'h0003,
16'h2D26, 16'h0003,
16'h2D27, 16'h0003,
16'h2D28, 16'h0003,
16'h2D29, 16'h0003,
16'h2D2A, 16'h0003,
16'h2D2B, 16'h0003,
16'h2D2C, 16'h0003,
16'h2D2D, 16'h0003,
16'h2D2E, 16'h0003,
16'h2D2F, 16'h0003,
16'h2D30, 16'h0003,
16'h2D31, 16'h0003,
16'h2D32, 16'h0003,
16'h2D33, 16'h0003,
16'h2D34, 16'h0003,
16'h2D35, 16'h0003,
16'h2D36, 16'h0003,
16'h2D37, 16'h0003,
16'h2D38, 16'h0003,
16'h2D39, 16'h0003,
16'h2D3A, 16'h0003,
16'h2D3B, 16'h0003,
16'h2D3C, 16'h0003,
16'h2D3D, 16'h0003,
16'h2D3E, 16'h0003,
16'h2D3F, 16'h0003,
16'h2D40, 16'h0003,
16'h2D41, 16'h0003,
16'h2D42, 16'h0003,
16'h2D43, 16'h0003,
16'h2D44, 16'h0003,
16'h2D45, 16'h0003,
16'h2D46, 16'h0003,
16'h2D47, 16'h0003,
16'h2D48, 16'h0003,
16'h2D49, 16'h0003,
16'h2D4A, 16'h0003,
16'h2D4B, 16'h0003,
16'h2D4C, 16'h0003,
16'h2D4D, 16'h0003,
16'h2D4E, 16'h0003,
16'h2D4F, 16'h0003,
16'h2D50, 16'h0003,
16'h2D51, 16'h0003,
16'h2D52, 16'h0003,
16'h2D53, 16'h0003,
16'h2D54, 16'h0003,
16'h2D55, 16'h0003,
16'h2D56, 16'h0003,
16'h2D57, 16'h0003,
16'h2D58, 16'h0003,
16'h2D59, 16'h0003,
16'h2D5A, 16'h0003,
16'h2D5B, 16'h0003,
16'h2D5C, 16'h0003,
16'h2D5D, 16'h0003,
16'h2D5E, 16'h0003,
16'h2D5F, 16'h0003,
16'h2D60, 16'h0003,
16'h2D61, 16'h0003,
16'h2D62, 16'h0003,
16'h2D63, 16'h0003,
16'h2D64, 16'h0003,
16'h2D65, 16'h0003,
16'h2D66, 16'h0003,
16'h2D67, 16'h0003,
16'h2D68, 16'h0003,
16'h2D69, 16'h0003,
16'h2D6A, 16'h0003,
16'h2D6B, 16'h0003,
16'h2D6C, 16'h0003,
16'h2D6D, 16'h0003,
16'h2D6E, 16'h0003,
16'h2D6F, 16'h0003,
16'h2D70, 16'h0003,
16'h2D71, 16'h0003,
16'h2D72, 16'h0003,
16'h2D73, 16'h0003,
16'h2D74, 16'h0003,
16'h2D75, 16'h0003,
16'h2D76, 16'h0003,
16'h2D77, 16'h0003,
16'h2D78, 16'h0003,
16'h2D79, 16'h0003,
16'h2D7A, 16'h0003,
16'h2D7B, 16'h0003,
16'h2D7C, 16'h0003,
16'h2D7D, 16'h0003,
16'h2D7E, 16'h0003,
16'h2D7F, 16'h0003,
16'h2D80, 16'h0003,
16'h2D81, 16'h0003,
16'h2D82, 16'h0003,
16'h2D83, 16'h0003,
16'h2D84, 16'h0003,
16'h2D85, 16'h0003,
16'h2D86, 16'h0003,
16'h2D87, 16'h0003,
16'h2D88, 16'h0003,
16'h2D89, 16'h0003,
16'h2D8A, 16'h0003,
16'h2D8B, 16'h0003,
16'h2D8C, 16'h0003,
16'h2D8D, 16'h0003,
16'h2D8E, 16'h0003,
16'h2D8F, 16'h0003,
16'h2D90, 16'h0003,
16'h2D91, 16'h0003,
16'h2D92, 16'h0003,
16'h2D93, 16'h0003,
16'h2D94, 16'h0003,
16'h2D95, 16'h0003,
16'h2D96, 16'h0003,
16'h2D97, 16'h0003,
16'h2D98, 16'h0003,
16'h2D99, 16'h0003,
16'h2D9A, 16'h0003,
16'h2D9B, 16'h0003,
16'h2D9C, 16'h0003,
16'h2D9D, 16'h0003,
16'h2D9E, 16'h0003,
16'h2D9F, 16'h0003,
16'h2DA0, 16'h0003,
16'h2DA1, 16'h0003,
16'h2DA2, 16'h0003,
16'h2DA3, 16'h0003,
16'h2DA4, 16'h0003,
16'h2DA5, 16'h0003,
16'h2DA6, 16'h0003,
16'h2DA7, 16'h0003,
16'h2DA8, 16'h0003,
16'h2DA9, 16'h0003,
16'h2DAA, 16'h0003,
16'h2DAB, 16'h0003,
16'h2DAC, 16'h0003,
16'h2DAD, 16'h0003,
16'h2DAE, 16'h0003,
16'h2DAF, 16'h0003,
16'h2DB0, 16'h0003,
16'h2DB1, 16'h0003,
16'h2DB2, 16'h0003,
16'h2DB3, 16'h0003,
16'h2DB4, 16'h0003,
16'h2DB5, 16'h0003,
16'h2DB6, 16'h0003,
16'h2DB7, 16'h0003,
16'h2DB8, 16'h0003,
16'h2DB9, 16'h0003,
16'h2DBA, 16'h0003,
16'h2DBB, 16'h0003,
16'h2DBC, 16'h0003,
16'h2DBD, 16'h0003,
16'h2DBE, 16'h0003,
16'h2DBF, 16'h0003,
16'h2DC0, 16'h0003,
16'h2DC1, 16'h0003,
16'h2DC2, 16'h0003,
16'h2DC3, 16'h0003,
16'h2DC4, 16'h0003,
16'h2DC5, 16'h0003,
16'h2DC6, 16'h0003,
16'h2DC7, 16'h0003,
16'h2DC8, 16'h0003,
16'h2DC9, 16'h0003,
16'h2DCA, 16'h0003,
16'h2DCB, 16'h0003,
16'h2DCC, 16'h0003,
16'h2DCD, 16'h0003,
16'h2DCE, 16'h0003,
16'h2DCF, 16'h0003,
16'h2DD0, 16'h0003,
16'h2DD1, 16'h0003,
16'h2DD2, 16'h0003,
16'h2DD3, 16'h0003,
16'h2DD4, 16'h0003,
16'h2DD5, 16'h0003,
16'h2DD6, 16'h0003,
16'h2DD7, 16'h0003,
16'h2DD8, 16'h0003,
16'h2DD9, 16'h0003,
16'h2DDA, 16'h0003,
16'h2DDB, 16'h0003,
16'h2DDC, 16'h0003,
16'h2DDD, 16'h0003,
16'h2DDE, 16'h0003,
16'h2DDF, 16'h0003,
16'h2DE0, 16'h0003,
16'h2DE1, 16'h0003,
16'h2DE2, 16'h0003,
16'h2DE3, 16'h0003,
16'h2DE4, 16'h0003,
16'h2DE5, 16'h0003,
16'h2DE6, 16'h0003,
16'h2DE7, 16'h0003,
16'h2DE8, 16'h0003,
16'h2DE9, 16'h0003,
16'h2DEA, 16'h0003,
16'h2DEB, 16'h0003,
16'h2DEC, 16'h0003,
16'h2DED, 16'h0003,
16'h2DEE, 16'h0003,
16'h2DEF, 16'h0003,
16'h2DF0, 16'h0003,
16'h2DF1, 16'h0003,
16'h2DF2, 16'h0003,
16'h2DF3, 16'h0003,
16'h2DF4, 16'h0003,
16'h2DF5, 16'h0003,
16'h2DF6, 16'h0003,
16'h2DF7, 16'h0003,
16'h2DF8, 16'h0003,
16'h2DF9, 16'h0003,
16'h2DFA, 16'h0003,
16'h2DFB, 16'h0003,
16'h2DFC, 16'h0003,
16'h2DFD, 16'h0003,
16'h2DFE, 16'h0003,
16'h2DFF, 16'h0003,
16'h2E00, 16'h0003,
16'h2E01, 16'h0003,
16'h2E02, 16'h0003,
16'h2E03, 16'h0003,
16'h2E04, 16'h0003,
16'h2E05, 16'h0003,
16'h2E06, 16'h0003,
16'h2E07, 16'h0003,
16'h2E08, 16'h0003,
16'h2E09, 16'h0003,
16'h2E0A, 16'h0003,
16'h2E0B, 16'h0003,
16'h2E0C, 16'h0003,
16'h2E0D, 16'h0003,
16'h2E0E, 16'h0003,
16'h2E0F, 16'h0003,
16'h2E10, 16'h0003,
16'h2E11, 16'h0003,
16'h2E12, 16'h0003,
16'h2E13, 16'h0003,
16'h2E14, 16'h0003,
16'h2E15, 16'h0003,
16'h2E16, 16'h0003,
16'h2E17, 16'h0003,
16'h2E18, 16'h0003,
16'h2E19, 16'h0003,
16'h2E1A, 16'h0003,
16'h2E1B, 16'h0003,
16'h2E1C, 16'h0003,
16'h2E1D, 16'h0003,
16'h2E1E, 16'h0003,
16'h2E1F, 16'h0003,
16'h2E20, 16'h0003,
16'h2E21, 16'h0003,
16'h2E22, 16'h0003,
16'h2E23, 16'h0003,
16'h2E24, 16'h0003,
16'h2E25, 16'h0003,
16'h2E26, 16'h0003,
16'h2E27, 16'h0003,
16'h2E28, 16'h0003,
16'h2E29, 16'h0003,
16'h2E2A, 16'h0003,
16'h2E2B, 16'h0003,
16'h2E2C, 16'h0003,
16'h2E2D, 16'h0003,
16'h2E2E, 16'h0003,
16'h2E2F, 16'h0003,
16'h2E30, 16'h0003,
16'h2E31, 16'h0003,
16'h2E32, 16'h0003,
16'h2E33, 16'h0003,
16'h2E34, 16'h0003,
16'h2E35, 16'h0003,
16'h2E36, 16'h0003,
16'h2E37, 16'h0003,
16'h2E38, 16'h0003,
16'h2E39, 16'h0003,
16'h2E3A, 16'h0003,
16'h2E3B, 16'h0003,
16'h2E3C, 16'h0003,
16'h2E3D, 16'h0003,
16'h2E3E, 16'h0003,
16'h2E3F, 16'h0003,
16'h2E40, 16'h0003,
16'h2E41, 16'h0003,
16'h2E42, 16'h0003,
16'h2E43, 16'h0003,
16'h2E44, 16'h0003,
16'h2E45, 16'h0003,
16'h2E46, 16'h0003,
16'h2E47, 16'h0003,
16'h2E48, 16'h0003,
16'h2E49, 16'h0003,
16'h2E4A, 16'h0003,
16'h2E4B, 16'h0003,
16'h2E4C, 16'h0003,
16'h2E4D, 16'h0003,
16'h2E4E, 16'h0003,
16'h2E4F, 16'h0003,
16'h2E50, 16'h0003,
16'h2E51, 16'h0003,
16'h2E52, 16'h0003,
16'h2E53, 16'h0003,
16'h2E54, 16'h0003,
16'h2E55, 16'h0003,
16'h2E56, 16'h0003,
16'h2E57, 16'h0003,
16'h2E58, 16'h0003,
16'h2E59, 16'h0003,
16'h2E5A, 16'h0003,
16'h2E5B, 16'h0003,
16'h2E5C, 16'h0003,
16'h2E5D, 16'h0003,
16'h2E5E, 16'h0003,
16'h2E5F, 16'h0003,
16'h2E60, 16'h0003,
16'h2E61, 16'h0003,
16'h2E62, 16'h0003,
16'h2E63, 16'h0003,
16'h2E64, 16'h0003,
16'h2E65, 16'h0003,
16'h2E66, 16'h0003,
16'h2E67, 16'h0003,
16'h2E68, 16'h0003,
16'h2E69, 16'h0003,
16'h2E6A, 16'h0003,
16'h2E6B, 16'h0003,
16'h2E6C, 16'h0003,
16'h2E6D, 16'h0003,
16'h2E6E, 16'h0003,
16'h2E6F, 16'h0003,
16'h2E70, 16'h0003,
16'h2E71, 16'h0003,
16'h2E72, 16'h0003,
16'h2E73, 16'h0003,
16'h2E74, 16'h0003,
16'h2E75, 16'h0003,
16'h2E76, 16'h0003,
16'h2E77, 16'h0003,
16'h2E78, 16'h0003,
16'h2E79, 16'h0003,
16'h2E7A, 16'h0003,
16'h2E7B, 16'h0003,
16'h2E7C, 16'h0003,
16'h2E7D, 16'h0003,
16'h2E7E, 16'h0003,
16'h2E7F, 16'h0003,
16'h2E80, 16'h0003,
16'h2E81, 16'h0003,
16'h2E82, 16'h0003,
16'h2E83, 16'h0003,
16'h2E84, 16'h0003,
16'h2E85, 16'h0003,
16'h2E86, 16'h0003,
16'h2E87, 16'h0003,
16'h2E88, 16'h0003,
16'h2E89, 16'h0003,
16'h2E8A, 16'h0003,
16'h2E8B, 16'h0003,
16'h2E8C, 16'h0003,
16'h2E8D, 16'h0003,
16'h2E8E, 16'h0003,
16'h2E8F, 16'h0003,
16'h2E90, 16'h0003,
16'h2E91, 16'h0003,
16'h2E92, 16'h0003,
16'h2E93, 16'h0003,
16'h2E94, 16'h0003,
16'h2E95, 16'h0003,
16'h2E96, 16'h0003,
16'h2E97, 16'h0003,
16'h2E98, 16'h0003,
16'h2E99, 16'h0003,
16'h2E9A, 16'h0003,
16'h2E9B, 16'h0003,
16'h2E9C, 16'h0003,
16'h2E9D, 16'h0003,
16'h2E9E, 16'h0003,
16'h2E9F, 16'h0003,
16'h2EA0, 16'h0003,
16'h2EA1, 16'h0003,
16'h2EA2, 16'h0003,
16'h2EA3, 16'h0003,
16'h2EA4, 16'h0003,
16'h2EA5, 16'h0003,
16'h2EA6, 16'h0003,
16'h2EA7, 16'h0003,
16'h2EA8, 16'h0003,
16'h2EA9, 16'h0003,
16'h2EAA, 16'h0003,
16'h2EAB, 16'h0003,
16'h2EAC, 16'h0003,
16'h2EAD, 16'h0003,
16'h2EAE, 16'h0003,
16'h2EAF, 16'h0003,
16'h2EB0, 16'h0003,
16'h2EB1, 16'h0003,
16'h2EB2, 16'h0003,
16'h2EB3, 16'h0003,
16'h2EB4, 16'h0003,
16'h2EB5, 16'h0003,
16'h2EB6, 16'h0003,
16'h2EB7, 16'h0003,
16'h2EB8, 16'h0003,
16'h2EB9, 16'h0003,
16'h2EBA, 16'h0003,
16'h2EBB, 16'h0003,
16'h2EBC, 16'h0003,
16'h2EBD, 16'h0003,
16'h2EBE, 16'h0003,
16'h2EBF, 16'h0003,
16'h2EC0, 16'h00FF,
16'h2EC1, 16'h00FF,
16'h2EC2, 16'h00FF,
16'h2EC3, 16'h00FF,
16'h2EC4, 16'h00FF,
16'h2EC5, 16'h00FF,
16'h2EC6, 16'h00FF,
16'h2EC7, 16'h00FF,
16'h2EC8, 16'h00FF,
16'h2EC9, 16'h00FF,
16'h2ECA, 16'h00FF,
16'h2ECB, 16'h00FF,
16'h2ECC, 16'h00FF,
16'h2ECD, 16'h00FF,
16'h2ECE, 16'h00FF,
16'h2ECF, 16'h00FF,
16'h2ED0, 16'h00FF,
16'h2ED1, 16'h00FF,
16'h2ED2, 16'h00FF,
16'h2ED3, 16'h00FF,
16'h2ED4, 16'h00FF,
16'h2ED5, 16'h00FF,
16'h2ED6, 16'h00FF,
16'h2ED7, 16'h00FF,
16'h2ED8, 16'h00FF,
16'h2ED9, 16'h00FF,
16'h2EDA, 16'h00FF,
16'h2EDB, 16'h00FF,
16'h2EDC, 16'h00FF,
16'h2EDD, 16'h00FF,
16'h2EDE, 16'h00FF,
16'h2EDF, 16'h00FF,
16'h2EE0, 16'h00FF,
16'h2EE1, 16'h00FF,
16'h2EE2, 16'h00FF,
16'h2EE3, 16'h00FF,
16'h2EE4, 16'h00FF,
16'h2EE5, 16'h00FF,
16'h2EE6, 16'h00FF,
16'h2EE7, 16'h00FF,
16'h2EE8, 16'h00FF,
16'h2EE9, 16'h00FF,
16'h2EEA, 16'h00FF,
16'h2EEB, 16'h00FF,
16'h2EEC, 16'h00FF,
16'h2EED, 16'h00FF,
16'h2EEE, 16'h00FF,
16'h2EEF, 16'h00FF,
16'h2EF0, 16'h00FF,
16'h2EF1, 16'h00FF,
16'h2EF2, 16'h00FF,
16'h2EF3, 16'h00FF,
16'h2EF4, 16'h00FF,
16'h2EF5, 16'h00FF,
16'h2EF6, 16'h00FF,
16'h2EF7, 16'h00FF,
16'h2EF8, 16'h00FF,
16'h2EF9, 16'h00FF,
16'h2EFA, 16'h00FF,
16'h2EFB, 16'h00FF,
16'h2EFC, 16'h00FF,
16'h2EFD, 16'h00FF,
16'h2EFE, 16'h00FF,
16'h2EFF, 16'h00FF,
16'h3F00, 16'h0000,
16'h3F01, 16'h0001,
16'h3F02, 16'h0002,
16'h3F03, 16'h0003,
16'h3F04, 16'h0004,
16'h3F05, 16'h0005,
16'h3F06, 16'h0006,
16'h3F07, 16'h0007,
16'h3F08, 16'h0008,
16'h3F09, 16'h0009,
16'h3F0A, 16'h000A,
16'h3F0B, 16'h000B,
16'h3F0C, 16'h000C,
16'h3F0D, 16'h000D,
16'h3F0E, 16'h000E,
16'h3F0F, 16'h000F,
16'h3F10, 16'h0010,
16'h3F11, 16'h0011,
16'h3F12, 16'h0012,
16'h3F13, 16'h0013,
16'h3F14, 16'h0014,
16'h3F15, 16'h0015,
16'h3F16, 16'h0016,
16'h3F17, 16'h0017,
16'h3F18, 16'h0018,
16'h3F19, 16'h0019,
16'h3F1A, 16'h001A,
16'h3F1B, 16'h001B,
16'h3F1C, 16'h001C,
16'h3F1D, 16'h001D,
16'h3F1E, 16'h001E,
16'h3F1F, 16'h001F



};


endpackage
