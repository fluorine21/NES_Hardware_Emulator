



module interrupt_handler_tb();





endmodule

