

package vram_listing;


integer spram_listing[64] = 
{
//Sprite 0
8'h00, 8'h00, //row 0
8'h01, 8'h00, // Tile 1F
8'h02, 8'h80, // Attribute bytes
8'h03, 8'h00, //Col 0

//Sprite 1
8'h04, 8'h08, //row 0
8'h05, 8'h00, // Tile 1F
8'h06, 8'h40, // Attribute bytes
8'h07, 8'h08, //Col 8

//Sprite 2
8'h08, 8'h10, //row 0
8'h09, 8'h00, // Tile 1F
8'h0A, 8'hC2, // Attribute bytes
8'h0B, 8'h10, //Col 16

//Sprite 3
8'h0C, 8'h18, //row 0
8'h0D, 8'h00, // Tile 1F
8'h0E, 8'h03, // Attribute bytes
8'h0F, 8'h18, //Col 24

//Sprite 4
8'h10, 8'h20, //row 0
8'h11, 8'h00, // Tile 1F
8'h12, 8'h00, // Attribute bytes
8'h13, 8'h20, //Col 32

//Sprite 5
8'h14, 8'h28, //row 0
8'h15, 8'h00, // Tile 1F
8'h16, 8'h01, // Attribute bytes
8'h17, 8'h28, //Col 40

//Sprite 6
8'h18, 8'h30, //row 0
8'h19, 8'h00, // Tile 1F
8'h1A, 8'h02, // Attribute bytes
8'h1B, 8'h30, //Col 48

//Sprite 7
8'h1C, 8'h38, //row 0
8'h1D, 8'h00, // Tile 1F
8'h1E, 8'h03, // Attribute bytes
8'h1F, 8'h38 //Col 56
};



integer vram_listing[] = 
{


16'h0000, 16'h0000,
16'h0001, 16'h00FF,
16'h0002, 16'h0000,
16'h0003, 16'h00FF,
16'h0004, 16'h0000,
16'h0005, 16'h00FF,
16'h0006, 16'h0000,
16'h0007, 16'h00FF,
16'h0008, 16'h0000,
16'h0009, 16'h00FF,
16'h000A, 16'h0000,
16'h000B, 16'h00FF,
16'h000C, 16'h0000,
16'h000D, 16'h00FF,
16'h000E, 16'h0000,
16'h000F, 16'h00FF,
16'h1000, 16'h0000,
16'h1001, 16'h00FF,
16'h1002, 16'h0000,
16'h1003, 16'h00FF,
16'h1004, 16'h0000,
16'h1005, 16'h00FF,
16'h1006, 16'h0000,
16'h1007, 16'h00FF,
16'h1008, 16'h0000,
16'h1009, 16'h00FF,
16'h100A, 16'h0000,
16'h100B, 16'h00FF,
16'h100C, 16'h0000,
16'h100D, 16'h00FF,
16'h100E, 16'h0000,
16'h100F, 16'h00FF,
16'h2000, 16'h0000,
16'h2001, 16'h0000,
16'h2002, 16'h0000,
16'h2003, 16'h0000,
16'h2004, 16'h0000,
16'h2005, 16'h0000,
16'h2006, 16'h0000,
16'h2007, 16'h0000,
16'h2008, 16'h0000,
16'h2009, 16'h0000,
16'h200A, 16'h0000,
16'h200B, 16'h0000,
16'h200C, 16'h0000,
16'h200D, 16'h0000,
16'h200E, 16'h0000,
16'h200F, 16'h0000,
16'h2010, 16'h0000,
16'h2011, 16'h0000,
16'h2012, 16'h0000,
16'h2013, 16'h0000,
16'h2014, 16'h0000,
16'h2015, 16'h0000,
16'h2016, 16'h0000,
16'h2017, 16'h0000,
16'h2018, 16'h0000,
16'h2019, 16'h0000,
16'h201A, 16'h0000,
16'h201B, 16'h0000,
16'h201C, 16'h0000,
16'h201D, 16'h0000,
16'h201E, 16'h0000,
16'h201F, 16'h0000,
16'h2020, 16'h0000,
16'h2021, 16'h0000,
16'h2022, 16'h0000,
16'h2023, 16'h0000,
16'h2024, 16'h0000,
16'h2025, 16'h0000,
16'h2026, 16'h0000,
16'h2027, 16'h0000,
16'h2028, 16'h0000,
16'h2029, 16'h0000,
16'h202A, 16'h0000,
16'h202B, 16'h0000,
16'h202C, 16'h0000,
16'h202D, 16'h0000,
16'h202E, 16'h0000,
16'h202F, 16'h0000,
16'h2030, 16'h0000,
16'h2031, 16'h0000,
16'h2032, 16'h0000,
16'h2033, 16'h0000,
16'h2034, 16'h0000,
16'h2035, 16'h0000,
16'h2036, 16'h0000,
16'h2037, 16'h0000,
16'h2038, 16'h0000,
16'h2039, 16'h0000,
16'h203A, 16'h0000,
16'h203B, 16'h0000,
16'h203C, 16'h0000,
16'h203D, 16'h0000,
16'h203E, 16'h0000,
16'h203F, 16'h0000,
16'h2040, 16'h0000,
16'h2041, 16'h0000,
16'h2042, 16'h0000,
16'h2043, 16'h0000,
16'h2044, 16'h0000,
16'h2045, 16'h0000,
16'h2046, 16'h0000,
16'h2047, 16'h0000,
16'h2048, 16'h0000,
16'h2049, 16'h0000,
16'h204A, 16'h0000,
16'h204B, 16'h0000,
16'h204C, 16'h0000,
16'h204D, 16'h0000,
16'h204E, 16'h0000,
16'h204F, 16'h0000,
16'h2050, 16'h0000,
16'h2051, 16'h0000,
16'h2052, 16'h0000,
16'h2053, 16'h0000,
16'h2054, 16'h0000,
16'h2055, 16'h0000,
16'h2056, 16'h0000,
16'h2057, 16'h0000,
16'h2058, 16'h0000,
16'h2059, 16'h0000,
16'h205A, 16'h0000,
16'h205B, 16'h0000,
16'h205C, 16'h0000,
16'h205D, 16'h0000,
16'h205E, 16'h0000,
16'h205F, 16'h0000,
16'h2060, 16'h0000,
16'h2061, 16'h0000,
16'h2062, 16'h0000,
16'h2063, 16'h0000,
16'h2064, 16'h0000,
16'h2065, 16'h0000,
16'h2066, 16'h0000,
16'h2067, 16'h0000,
16'h2068, 16'h0000,
16'h2069, 16'h0000,
16'h206A, 16'h0000,
16'h206B, 16'h0000,
16'h206C, 16'h0000,
16'h206D, 16'h0000,
16'h206E, 16'h0000,
16'h206F, 16'h0000,
16'h2070, 16'h0000,
16'h2071, 16'h0000,
16'h2072, 16'h0000,
16'h2073, 16'h0000,
16'h2074, 16'h0000,
16'h2075, 16'h0000,
16'h2076, 16'h0000,
16'h2077, 16'h0000,
16'h2078, 16'h0000,
16'h2079, 16'h0000,
16'h207A, 16'h0000,
16'h207B, 16'h0000,
16'h207C, 16'h0000,
16'h207D, 16'h0000,
16'h207E, 16'h0000,
16'h207F, 16'h0000,
16'h2080, 16'h0000,
16'h2081, 16'h0000,
16'h2082, 16'h0000,
16'h2083, 16'h0000,
16'h2084, 16'h0000,
16'h2085, 16'h0000,
16'h2086, 16'h0000,
16'h2087, 16'h0000,
16'h2088, 16'h0000,
16'h2089, 16'h0000,
16'h208A, 16'h0000,
16'h208B, 16'h0000,
16'h208C, 16'h0000,
16'h208D, 16'h0000,
16'h208E, 16'h0000,
16'h208F, 16'h0000,
16'h2090, 16'h0000,
16'h2091, 16'h0000,
16'h2092, 16'h0000,
16'h2093, 16'h0000,
16'h2094, 16'h0000,
16'h2095, 16'h0000,
16'h2096, 16'h0000,
16'h2097, 16'h0000,
16'h2098, 16'h0000,
16'h2099, 16'h0000,
16'h209A, 16'h0000,
16'h209B, 16'h0000,
16'h209C, 16'h0000,
16'h209D, 16'h0000,
16'h209E, 16'h0000,
16'h209F, 16'h0000,
16'h20A0, 16'h0000,
16'h20A1, 16'h0000,
16'h20A2, 16'h0000,
16'h20A3, 16'h0000,
16'h20A4, 16'h0000,
16'h20A5, 16'h0000,
16'h20A6, 16'h0000,
16'h20A7, 16'h0000,
16'h20A8, 16'h0000,
16'h20A9, 16'h0000,
16'h20AA, 16'h0000,
16'h20AB, 16'h0000,
16'h20AC, 16'h0000,
16'h20AD, 16'h0000,
16'h20AE, 16'h0000,
16'h20AF, 16'h0000,
16'h20B0, 16'h0000,
16'h20B1, 16'h0000,
16'h20B2, 16'h0000,
16'h20B3, 16'h0000,
16'h20B4, 16'h0000,
16'h20B5, 16'h0000,
16'h20B6, 16'h0000,
16'h20B7, 16'h0000,
16'h20B8, 16'h0000,
16'h20B9, 16'h0000,
16'h20BA, 16'h0000,
16'h20BB, 16'h0000,
16'h20BC, 16'h0000,
16'h20BD, 16'h0000,
16'h20BE, 16'h0000,
16'h20BF, 16'h0000,
16'h20C0, 16'h0000,
16'h20C1, 16'h0000,
16'h20C2, 16'h0000,
16'h20C3, 16'h0000,
16'h20C4, 16'h0000,
16'h20C5, 16'h0000,
16'h20C6, 16'h0000,
16'h20C7, 16'h0000,
16'h20C8, 16'h0000,
16'h20C9, 16'h0000,
16'h20CA, 16'h0000,
16'h20CB, 16'h0000,
16'h20CC, 16'h0000,
16'h20CD, 16'h0000,
16'h20CE, 16'h0000,
16'h20CF, 16'h0000,
16'h20D0, 16'h0000,
16'h20D1, 16'h0000,
16'h20D2, 16'h0000,
16'h20D3, 16'h0000,
16'h20D4, 16'h0000,
16'h20D5, 16'h0000,
16'h20D6, 16'h0000,
16'h20D7, 16'h0000,
16'h20D8, 16'h0000,
16'h20D9, 16'h0000,
16'h20DA, 16'h0000,
16'h20DB, 16'h0000,
16'h20DC, 16'h0000,
16'h20DD, 16'h0000,
16'h20DE, 16'h0000,
16'h20DF, 16'h0000,
16'h20E0, 16'h0000,
16'h20E1, 16'h0000,
16'h20E2, 16'h0000,
16'h20E3, 16'h0000,
16'h20E4, 16'h0000,
16'h20E5, 16'h0000,
16'h20E6, 16'h0000,
16'h20E7, 16'h0000,
16'h20E8, 16'h0000,
16'h20E9, 16'h0000,
16'h20EA, 16'h0000,
16'h20EB, 16'h0000,
16'h20EC, 16'h0000,
16'h20ED, 16'h0000,
16'h20EE, 16'h0000,
16'h20EF, 16'h0000,
16'h20F0, 16'h0000,
16'h20F1, 16'h0000,
16'h20F2, 16'h0000,
16'h20F3, 16'h0000,
16'h20F4, 16'h0000,
16'h20F5, 16'h0000,
16'h20F6, 16'h0000,
16'h20F7, 16'h0000,
16'h20F8, 16'h0000,
16'h20F9, 16'h0000,
16'h20FA, 16'h0000,
16'h20FB, 16'h0000,
16'h20FC, 16'h0000,
16'h20FD, 16'h0000,
16'h20FE, 16'h0000,
16'h20FF, 16'h0000,
16'h2100, 16'h0000,
16'h2101, 16'h0000,
16'h2102, 16'h0000,
16'h2103, 16'h0000,
16'h2104, 16'h0000,
16'h2105, 16'h0000,
16'h2106, 16'h0000,
16'h2107, 16'h0000,
16'h2108, 16'h0000,
16'h2109, 16'h0000,
16'h210A, 16'h0000,
16'h210B, 16'h0000,
16'h210C, 16'h0000,
16'h210D, 16'h0000,
16'h210E, 16'h0000,
16'h210F, 16'h0000,
16'h2110, 16'h0000,
16'h2111, 16'h0000,
16'h2112, 16'h0000,
16'h2113, 16'h0000,
16'h2114, 16'h0000,
16'h2115, 16'h0000,
16'h2116, 16'h0000,
16'h2117, 16'h0000,
16'h2118, 16'h0000,
16'h2119, 16'h0000,
16'h211A, 16'h0000,
16'h211B, 16'h0000,
16'h211C, 16'h0000,
16'h211D, 16'h0000,
16'h211E, 16'h0000,
16'h211F, 16'h0000,
16'h2120, 16'h0000,
16'h2121, 16'h0000,
16'h2122, 16'h0000,
16'h2123, 16'h0000,
16'h2124, 16'h0000,
16'h2125, 16'h0000,
16'h2126, 16'h0000,
16'h2127, 16'h0000,
16'h2128, 16'h0000,
16'h2129, 16'h0000,
16'h212A, 16'h0000,
16'h212B, 16'h0000,
16'h212C, 16'h0000,
16'h212D, 16'h0000,
16'h212E, 16'h0000,
16'h212F, 16'h0000,
16'h2130, 16'h0000,
16'h2131, 16'h0000,
16'h2132, 16'h0000,
16'h2133, 16'h0000,
16'h2134, 16'h0000,
16'h2135, 16'h0000,
16'h2136, 16'h0000,
16'h2137, 16'h0000,
16'h2138, 16'h0000,
16'h2139, 16'h0000,
16'h213A, 16'h0000,
16'h213B, 16'h0000,
16'h213C, 16'h0000,
16'h213D, 16'h0000,
16'h213E, 16'h0000,
16'h213F, 16'h0000,
16'h2140, 16'h0000,
16'h2141, 16'h0000,
16'h2142, 16'h0000,
16'h2143, 16'h0000,
16'h2144, 16'h0000,
16'h2145, 16'h0000,
16'h2146, 16'h0000,
16'h2147, 16'h0000,
16'h2148, 16'h0000,
16'h2149, 16'h0000,
16'h214A, 16'h0000,
16'h214B, 16'h0000,
16'h214C, 16'h0000,
16'h214D, 16'h0000,
16'h214E, 16'h0000,
16'h214F, 16'h0000,
16'h2150, 16'h0000,
16'h2151, 16'h0000,
16'h2152, 16'h0000,
16'h2153, 16'h0000,
16'h2154, 16'h0000,
16'h2155, 16'h0000,
16'h2156, 16'h0000,
16'h2157, 16'h0000,
16'h2158, 16'h0000,
16'h2159, 16'h0000,
16'h215A, 16'h0000,
16'h215B, 16'h0000,
16'h215C, 16'h0000,
16'h215D, 16'h0000,
16'h215E, 16'h0000,
16'h215F, 16'h0000,
16'h2160, 16'h0000,
16'h2161, 16'h0000,
16'h2162, 16'h0000,
16'h2163, 16'h0000,
16'h2164, 16'h0000,
16'h2165, 16'h0000,
16'h2166, 16'h0000,
16'h2167, 16'h0000,
16'h2168, 16'h0000,
16'h2169, 16'h0000,
16'h216A, 16'h0000,
16'h216B, 16'h0000,
16'h216C, 16'h0000,
16'h216D, 16'h0000,
16'h216E, 16'h0000,
16'h216F, 16'h0000,
16'h2170, 16'h0000,
16'h2171, 16'h0000,
16'h2172, 16'h0000,
16'h2173, 16'h0000,
16'h2174, 16'h0000,
16'h2175, 16'h0000,
16'h2176, 16'h0000,
16'h2177, 16'h0000,
16'h2178, 16'h0000,
16'h2179, 16'h0000,
16'h217A, 16'h0000,
16'h217B, 16'h0000,
16'h217C, 16'h0000,
16'h217D, 16'h0000,
16'h217E, 16'h0000,
16'h217F, 16'h0000,
16'h2180, 16'h0000,
16'h2181, 16'h0000,
16'h2182, 16'h0000,
16'h2183, 16'h0000,
16'h2184, 16'h0000,
16'h2185, 16'h0000,
16'h2186, 16'h0000,
16'h2187, 16'h0000,
16'h2188, 16'h0000,
16'h2189, 16'h0000,
16'h218A, 16'h0000,
16'h218B, 16'h0000,
16'h218C, 16'h0000,
16'h218D, 16'h0000,
16'h218E, 16'h0000,
16'h218F, 16'h0000,
16'h2190, 16'h0000,
16'h2191, 16'h0000,
16'h2192, 16'h0000,
16'h2193, 16'h0000,
16'h2194, 16'h0000,
16'h2195, 16'h0000,
16'h2196, 16'h0000,
16'h2197, 16'h0000,
16'h2198, 16'h0000,
16'h2199, 16'h0000,
16'h219A, 16'h0000,
16'h219B, 16'h0000,
16'h219C, 16'h0000,
16'h219D, 16'h0000,
16'h219E, 16'h0000,
16'h219F, 16'h0000,
16'h21A0, 16'h0000,
16'h21A1, 16'h0000,
16'h21A2, 16'h0000,
16'h21A3, 16'h0000,
16'h21A4, 16'h0000,
16'h21A5, 16'h0000,
16'h21A6, 16'h0000,
16'h21A7, 16'h0000,
16'h21A8, 16'h0000,
16'h21A9, 16'h0000,
16'h21AA, 16'h0000,
16'h21AB, 16'h0000,
16'h21AC, 16'h0000,
16'h21AD, 16'h0000,
16'h21AE, 16'h0000,
16'h21AF, 16'h0000,
16'h21B0, 16'h0000,
16'h21B1, 16'h0000,
16'h21B2, 16'h0000,
16'h21B3, 16'h0000,
16'h21B4, 16'h0000,
16'h21B5, 16'h0000,
16'h21B6, 16'h0000,
16'h21B7, 16'h0000,
16'h21B8, 16'h0000,
16'h21B9, 16'h0000,
16'h21BA, 16'h0000,
16'h21BB, 16'h0000,
16'h21BC, 16'h0000,
16'h21BD, 16'h0000,
16'h21BE, 16'h0000,
16'h21BF, 16'h0000,
16'h21C0, 16'h0000,
16'h21C1, 16'h0000,
16'h21C2, 16'h0000,
16'h21C3, 16'h0000,
16'h21C4, 16'h0000,
16'h21C5, 16'h0000,
16'h21C6, 16'h0000,
16'h21C7, 16'h0000,
16'h21C8, 16'h0000,
16'h21C9, 16'h0000,
16'h21CA, 16'h0000,
16'h21CB, 16'h0000,
16'h21CC, 16'h0000,
16'h21CD, 16'h0000,
16'h21CE, 16'h0000,
16'h21CF, 16'h0000,
16'h21D0, 16'h0000,
16'h21D1, 16'h0000,
16'h21D2, 16'h0000,
16'h21D3, 16'h0000,
16'h21D4, 16'h0000,
16'h21D5, 16'h0000,
16'h21D6, 16'h0000,
16'h21D7, 16'h0000,
16'h21D8, 16'h0000,
16'h21D9, 16'h0000,
16'h21DA, 16'h0000,
16'h21DB, 16'h0000,
16'h21DC, 16'h0000,
16'h21DD, 16'h0000,
16'h21DE, 16'h0000,
16'h21DF, 16'h0000,
16'h21E0, 16'h0000,
16'h21E1, 16'h0000,
16'h21E2, 16'h0000,
16'h21E3, 16'h0000,
16'h21E4, 16'h0000,
16'h21E5, 16'h0000,
16'h21E6, 16'h0000,
16'h21E7, 16'h0000,
16'h21E8, 16'h0000,
16'h21E9, 16'h0000,
16'h21EA, 16'h0000,
16'h21EB, 16'h0000,
16'h21EC, 16'h0000,
16'h21ED, 16'h0000,
16'h21EE, 16'h0000,
16'h21EF, 16'h0000,
16'h21F0, 16'h0000,
16'h21F1, 16'h0000,
16'h21F2, 16'h0000,
16'h21F3, 16'h0000,
16'h21F4, 16'h0000,
16'h21F5, 16'h0000,
16'h21F6, 16'h0000,
16'h21F7, 16'h0000,
16'h21F8, 16'h0000,
16'h21F9, 16'h0000,
16'h21FA, 16'h0000,
16'h21FB, 16'h0000,
16'h21FC, 16'h0000,
16'h21FD, 16'h0000,
16'h21FE, 16'h0000,
16'h21FF, 16'h0000,
16'h2200, 16'h0000,
16'h2201, 16'h0000,
16'h2202, 16'h0000,
16'h2203, 16'h0000,
16'h2204, 16'h0000,
16'h2205, 16'h0000,
16'h2206, 16'h0000,
16'h2207, 16'h0000,
16'h2208, 16'h0000,
16'h2209, 16'h0000,
16'h220A, 16'h0000,
16'h220B, 16'h0000,
16'h220C, 16'h0000,
16'h220D, 16'h0000,
16'h220E, 16'h0000,
16'h220F, 16'h0000,
16'h2210, 16'h0000,
16'h2211, 16'h0000,
16'h2212, 16'h0000,
16'h2213, 16'h0000,
16'h2214, 16'h0000,
16'h2215, 16'h0000,
16'h2216, 16'h0000,
16'h2217, 16'h0000,
16'h2218, 16'h0000,
16'h2219, 16'h0000,
16'h221A, 16'h0000,
16'h221B, 16'h0000,
16'h221C, 16'h0000,
16'h221D, 16'h0000,
16'h221E, 16'h0000,
16'h221F, 16'h0000,
16'h2220, 16'h0000,
16'h2221, 16'h0000,
16'h2222, 16'h0000,
16'h2223, 16'h0000,
16'h2224, 16'h0000,
16'h2225, 16'h0000,
16'h2226, 16'h0000,
16'h2227, 16'h0000,
16'h2228, 16'h0000,
16'h2229, 16'h0000,
16'h222A, 16'h0000,
16'h222B, 16'h0000,
16'h222C, 16'h0000,
16'h222D, 16'h0000,
16'h222E, 16'h0000,
16'h222F, 16'h0000,
16'h2230, 16'h0000,
16'h2231, 16'h0000,
16'h2232, 16'h0000,
16'h2233, 16'h0000,
16'h2234, 16'h0000,
16'h2235, 16'h0000,
16'h2236, 16'h0000,
16'h2237, 16'h0000,
16'h2238, 16'h0000,
16'h2239, 16'h0000,
16'h223A, 16'h0000,
16'h223B, 16'h0000,
16'h223C, 16'h0000,
16'h223D, 16'h0000,
16'h223E, 16'h0000,
16'h223F, 16'h0000,
16'h2240, 16'h0000,
16'h2241, 16'h0000,
16'h2242, 16'h0000,
16'h2243, 16'h0000,
16'h2244, 16'h0000,
16'h2245, 16'h0000,
16'h2246, 16'h0000,
16'h2247, 16'h0000,
16'h2248, 16'h0000,
16'h2249, 16'h0000,
16'h224A, 16'h0000,
16'h224B, 16'h0000,
16'h224C, 16'h0000,
16'h224D, 16'h0000,
16'h224E, 16'h0000,
16'h224F, 16'h0000,
16'h2250, 16'h0000,
16'h2251, 16'h0000,
16'h2252, 16'h0000,
16'h2253, 16'h0000,
16'h2254, 16'h0000,
16'h2255, 16'h0000,
16'h2256, 16'h0000,
16'h2257, 16'h0000,
16'h2258, 16'h0000,
16'h2259, 16'h0000,
16'h225A, 16'h0000,
16'h225B, 16'h0000,
16'h225C, 16'h0000,
16'h225D, 16'h0000,
16'h225E, 16'h0000,
16'h225F, 16'h0000,
16'h2260, 16'h0000,
16'h2261, 16'h0000,
16'h2262, 16'h0000,
16'h2263, 16'h0000,
16'h2264, 16'h0000,
16'h2265, 16'h0000,
16'h2266, 16'h0000,
16'h2267, 16'h0000,
16'h2268, 16'h0000,
16'h2269, 16'h0000,
16'h226A, 16'h0000,
16'h226B, 16'h0000,
16'h226C, 16'h0000,
16'h226D, 16'h0000,
16'h226E, 16'h0000,
16'h226F, 16'h0000,
16'h2270, 16'h0000,
16'h2271, 16'h0000,
16'h2272, 16'h0000,
16'h2273, 16'h0000,
16'h2274, 16'h0000,
16'h2275, 16'h0000,
16'h2276, 16'h0000,
16'h2277, 16'h0000,
16'h2278, 16'h0000,
16'h2279, 16'h0000,
16'h227A, 16'h0000,
16'h227B, 16'h0000,
16'h227C, 16'h0000,
16'h227D, 16'h0000,
16'h227E, 16'h0000,
16'h227F, 16'h0000,
16'h2280, 16'h0000,
16'h2281, 16'h0000,
16'h2282, 16'h0000,
16'h2283, 16'h0000,
16'h2284, 16'h0000,
16'h2285, 16'h0000,
16'h2286, 16'h0000,
16'h2287, 16'h0000,
16'h2288, 16'h0000,
16'h2289, 16'h0000,
16'h228A, 16'h0000,
16'h228B, 16'h0000,
16'h228C, 16'h0000,
16'h228D, 16'h0000,
16'h228E, 16'h0000,
16'h228F, 16'h0000,
16'h2290, 16'h0000,
16'h2291, 16'h0000,
16'h2292, 16'h0000,
16'h2293, 16'h0000,
16'h2294, 16'h0000,
16'h2295, 16'h0000,
16'h2296, 16'h0000,
16'h2297, 16'h0000,
16'h2298, 16'h0000,
16'h2299, 16'h0000,
16'h229A, 16'h0000,
16'h229B, 16'h0000,
16'h229C, 16'h0000,
16'h229D, 16'h0000,
16'h229E, 16'h0000,
16'h229F, 16'h0000,
16'h22A0, 16'h0000,
16'h22A1, 16'h0000,
16'h22A2, 16'h0000,
16'h22A3, 16'h0000,
16'h22A4, 16'h0000,
16'h22A5, 16'h0000,
16'h22A6, 16'h0000,
16'h22A7, 16'h0000,
16'h22A8, 16'h0000,
16'h22A9, 16'h0000,
16'h22AA, 16'h0000,
16'h22AB, 16'h0000,
16'h22AC, 16'h0000,
16'h22AD, 16'h0000,
16'h22AE, 16'h0000,
16'h22AF, 16'h0000,
16'h22B0, 16'h0000,
16'h22B1, 16'h0000,
16'h22B2, 16'h0000,
16'h22B3, 16'h0000,
16'h22B4, 16'h0000,
16'h22B5, 16'h0000,
16'h22B6, 16'h0000,
16'h22B7, 16'h0000,
16'h22B8, 16'h0000,
16'h22B9, 16'h0000,
16'h22BA, 16'h0000,
16'h22BB, 16'h0000,
16'h22BC, 16'h0000,
16'h22BD, 16'h0000,
16'h22BE, 16'h0000,
16'h22BF, 16'h0000,
16'h22C0, 16'h0000,
16'h22C1, 16'h0000,
16'h22C2, 16'h0000,
16'h22C3, 16'h0000,
16'h22C4, 16'h0000,
16'h22C5, 16'h0000,
16'h22C6, 16'h0000,
16'h22C7, 16'h0000,
16'h22C8, 16'h0000,
16'h22C9, 16'h0000,
16'h22CA, 16'h0000,
16'h22CB, 16'h0000,
16'h22CC, 16'h0000,
16'h22CD, 16'h0000,
16'h22CE, 16'h0000,
16'h22CF, 16'h0000,
16'h22D0, 16'h0000,
16'h22D1, 16'h0000,
16'h22D2, 16'h0000,
16'h22D3, 16'h0000,
16'h22D4, 16'h0000,
16'h22D5, 16'h0000,
16'h22D6, 16'h0000,
16'h22D7, 16'h0000,
16'h22D8, 16'h0000,
16'h22D9, 16'h0000,
16'h22DA, 16'h0000,
16'h22DB, 16'h0000,
16'h22DC, 16'h0000,
16'h22DD, 16'h0000,
16'h22DE, 16'h0000,
16'h22DF, 16'h0000,
16'h22E0, 16'h0000,
16'h22E1, 16'h0000,
16'h22E2, 16'h0000,
16'h22E3, 16'h0000,
16'h22E4, 16'h0000,
16'h22E5, 16'h0000,
16'h22E6, 16'h0000,
16'h22E7, 16'h0000,
16'h22E8, 16'h0000,
16'h22E9, 16'h0000,
16'h22EA, 16'h0000,
16'h22EB, 16'h0000,
16'h22EC, 16'h0000,
16'h22ED, 16'h0000,
16'h22EE, 16'h0000,
16'h22EF, 16'h0000,
16'h22F0, 16'h0000,
16'h22F1, 16'h0000,
16'h22F2, 16'h0000,
16'h22F3, 16'h0000,
16'h22F4, 16'h0000,
16'h22F5, 16'h0000,
16'h22F6, 16'h0000,
16'h22F7, 16'h0000,
16'h22F8, 16'h0000,
16'h22F9, 16'h0000,
16'h22FA, 16'h0000,
16'h22FB, 16'h0000,
16'h22FC, 16'h0000,
16'h22FD, 16'h0000,
16'h22FE, 16'h0000,
16'h22FF, 16'h0000,
16'h2300, 16'h0000,
16'h2301, 16'h0000,
16'h2302, 16'h0000,
16'h2303, 16'h0000,
16'h2304, 16'h0000,
16'h2305, 16'h0000,
16'h2306, 16'h0000,
16'h2307, 16'h0000,
16'h2308, 16'h0000,
16'h2309, 16'h0000,
16'h230A, 16'h0000,
16'h230B, 16'h0000,
16'h230C, 16'h0000,
16'h230D, 16'h0000,
16'h230E, 16'h0000,
16'h230F, 16'h0000,
16'h2310, 16'h0000,
16'h2311, 16'h0000,
16'h2312, 16'h0000,
16'h2313, 16'h0000,
16'h2314, 16'h0000,
16'h2315, 16'h0000,
16'h2316, 16'h0000,
16'h2317, 16'h0000,
16'h2318, 16'h0000,
16'h2319, 16'h0000,
16'h231A, 16'h0000,
16'h231B, 16'h0000,
16'h231C, 16'h0000,
16'h231D, 16'h0000,
16'h231E, 16'h0000,
16'h231F, 16'h0000,
16'h2320, 16'h0000,
16'h2321, 16'h0000,
16'h2322, 16'h0000,
16'h2323, 16'h0000,
16'h2324, 16'h0000,
16'h2325, 16'h0000,
16'h2326, 16'h0000,
16'h2327, 16'h0000,
16'h2328, 16'h0000,
16'h2329, 16'h0000,
16'h232A, 16'h0000,
16'h232B, 16'h0000,
16'h232C, 16'h0000,
16'h232D, 16'h0000,
16'h232E, 16'h0000,
16'h232F, 16'h0000,
16'h2330, 16'h0000,
16'h2331, 16'h0000,
16'h2332, 16'h0000,
16'h2333, 16'h0000,
16'h2334, 16'h0000,
16'h2335, 16'h0000,
16'h2336, 16'h0000,
16'h2337, 16'h0000,
16'h2338, 16'h0000,
16'h2339, 16'h0000,
16'h233A, 16'h0000,
16'h233B, 16'h0000,
16'h233C, 16'h0000,
16'h233D, 16'h0000,
16'h233E, 16'h0000,
16'h233F, 16'h0000,
16'h2340, 16'h0000,
16'h2341, 16'h0000,
16'h2342, 16'h0000,
16'h2343, 16'h0000,
16'h2344, 16'h0000,
16'h2345, 16'h0000,
16'h2346, 16'h0000,
16'h2347, 16'h0000,
16'h2348, 16'h0000,
16'h2349, 16'h0000,
16'h234A, 16'h0000,
16'h234B, 16'h0000,
16'h234C, 16'h0000,
16'h234D, 16'h0000,
16'h234E, 16'h0000,
16'h234F, 16'h0000,
16'h2350, 16'h0000,
16'h2351, 16'h0000,
16'h2352, 16'h0000,
16'h2353, 16'h0000,
16'h2354, 16'h0000,
16'h2355, 16'h0000,
16'h2356, 16'h0000,
16'h2357, 16'h0000,
16'h2358, 16'h0000,
16'h2359, 16'h0000,
16'h235A, 16'h0000,
16'h235B, 16'h0000,
16'h235C, 16'h0000,
16'h235D, 16'h0000,
16'h235E, 16'h0000,
16'h235F, 16'h0000,
16'h2360, 16'h0000,
16'h2361, 16'h0000,
16'h2362, 16'h0000,
16'h2363, 16'h0000,
16'h2364, 16'h0000,
16'h2365, 16'h0000,
16'h2366, 16'h0000,
16'h2367, 16'h0000,
16'h2368, 16'h0000,
16'h2369, 16'h0000,
16'h236A, 16'h0000,
16'h236B, 16'h0000,
16'h236C, 16'h0000,
16'h236D, 16'h0000,
16'h236E, 16'h0000,
16'h236F, 16'h0000,
16'h2370, 16'h0000,
16'h2371, 16'h0000,
16'h2372, 16'h0000,
16'h2373, 16'h0000,
16'h2374, 16'h0000,
16'h2375, 16'h0000,
16'h2376, 16'h0000,
16'h2377, 16'h0000,
16'h2378, 16'h0000,
16'h2379, 16'h0000,
16'h237A, 16'h0000,
16'h237B, 16'h0000,
16'h237C, 16'h0000,
16'h237D, 16'h0000,
16'h237E, 16'h0000,
16'h237F, 16'h0000,
16'h2380, 16'h0000,
16'h2381, 16'h0000,
16'h2382, 16'h0000,
16'h2383, 16'h0000,
16'h2384, 16'h0000,
16'h2385, 16'h0000,
16'h2386, 16'h0000,
16'h2387, 16'h0000,
16'h2388, 16'h0000,
16'h2389, 16'h0000,
16'h238A, 16'h0000,
16'h238B, 16'h0000,
16'h238C, 16'h0000,
16'h238D, 16'h0000,
16'h238E, 16'h0000,
16'h238F, 16'h0000,
16'h2390, 16'h0000,
16'h2391, 16'h0000,
16'h2392, 16'h0000,
16'h2393, 16'h0000,
16'h2394, 16'h0000,
16'h2395, 16'h0000,
16'h2396, 16'h0000,
16'h2397, 16'h0000,
16'h2398, 16'h0000,
16'h2399, 16'h0000,
16'h239A, 16'h0000,
16'h239B, 16'h0000,
16'h239C, 16'h0000,
16'h239D, 16'h0000,
16'h239E, 16'h0000,
16'h239F, 16'h0000,
16'h23A0, 16'h0000,
16'h23A1, 16'h0000,
16'h23A2, 16'h0000,
16'h23A3, 16'h0000,
16'h23A4, 16'h0000,
16'h23A5, 16'h0000,
16'h23A6, 16'h0000,
16'h23A7, 16'h0000,
16'h23A8, 16'h0000,
16'h23A9, 16'h0000,
16'h23AA, 16'h0000,
16'h23AB, 16'h0000,
16'h23AC, 16'h0000,
16'h23AD, 16'h0000,
16'h23AE, 16'h0000,
16'h23AF, 16'h0000,
16'h23B0, 16'h0000,
16'h23B1, 16'h0000,
16'h23B2, 16'h0000,
16'h23B3, 16'h0000,
16'h23B4, 16'h0000,
16'h23B5, 16'h0000,
16'h23B6, 16'h0000,
16'h23B7, 16'h0000,
16'h23B8, 16'h0000,
16'h23B9, 16'h0000,
16'h23BA, 16'h0000,
16'h23BB, 16'h0000,
16'h23BC, 16'h0000,
16'h23BD, 16'h0000,
16'h23BE, 16'h0000,
16'h23BF, 16'h0000,
16'h23C0, 16'h0000,
16'h23C1, 16'h0000,
16'h23C2, 16'h0000,
16'h23C3, 16'h0000,
16'h23C4, 16'h0000,
16'h23C5, 16'h0000,
16'h23C6, 16'h0000,
16'h23C7, 16'h0000,
16'h23C8, 16'h0000,
16'h23C9, 16'h0000,
16'h23CA, 16'h0000,
16'h23CB, 16'h0000,
16'h23CC, 16'h0000,
16'h23CD, 16'h0000,
16'h23CE, 16'h0000,
16'h23CF, 16'h0000,
16'h23D0, 16'h0000,
16'h23D1, 16'h0000,
16'h23D2, 16'h0000,
16'h23D3, 16'h0000,
16'h23D4, 16'h0000,
16'h23D5, 16'h0000,
16'h23D6, 16'h0000,
16'h23D7, 16'h0000,
16'h23D8, 16'h0000,
16'h23D9, 16'h0000,
16'h23DA, 16'h0000,
16'h23DB, 16'h0000,
16'h23DC, 16'h0000,
16'h23DD, 16'h0000,
16'h23DE, 16'h0000,
16'h23DF, 16'h0000,
16'h23E0, 16'h0000,
16'h23E1, 16'h0000,
16'h23E2, 16'h0000,
16'h23E3, 16'h0000,
16'h23E4, 16'h0000,
16'h23E5, 16'h0000,
16'h23E6, 16'h0000,
16'h23E7, 16'h0000,
16'h23E8, 16'h0000,
16'h23E9, 16'h0000,
16'h23EA, 16'h0000,
16'h23EB, 16'h0000,
16'h23EC, 16'h0000,
16'h23ED, 16'h0000,
16'h23EE, 16'h0000,
16'h23EF, 16'h0000,
16'h23F0, 16'h0000,
16'h23F1, 16'h0000,
16'h23F2, 16'h0000,
16'h23F3, 16'h0000,
16'h23F4, 16'h0000,
16'h23F5, 16'h0000,
16'h23F6, 16'h0000,
16'h23F7, 16'h0000,
16'h23F8, 16'h0000,
16'h23F9, 16'h0000,
16'h23FA, 16'h0000,
16'h23FB, 16'h0000,
16'h23FC, 16'h0000,
16'h23FD, 16'h0000,
16'h23FE, 16'h0000,
16'h23FF, 16'h0000,
16'h3F00, 16'h0000,
16'h3F01, 16'h0001,
16'h3F02, 16'h0002,
16'h3F03, 16'h0003,
16'h3F04, 16'h0004,
16'h3F05, 16'h0005,
16'h3F06, 16'h0006,
16'h3F07, 16'h0007,
16'h3F08, 16'h0008,
16'h3F09, 16'h0009,
16'h3F0A, 16'h000A,
16'h3F0B, 16'h000B,
16'h3F0C, 16'h000C,
16'h3F0D, 16'h000D,
16'h3F0E, 16'h000E,
16'h3F0F, 16'h000F,
16'h3F10, 16'h0010,
16'h3F11, 16'h0011,
16'h3F12, 16'h0012,
16'h3F13, 16'h0013,
16'h3F14, 16'h0014,
16'h3F15, 16'h0015,
16'h3F16, 16'h0016,
16'h3F17, 16'h0017,
16'h3F18, 16'h0018,
16'h3F19, 16'h0019,
16'h3F1A, 16'h001A,
16'h3F1B, 16'h001B,
16'h3F1C, 16'h001C,
16'h3F1D, 16'h001D,
16'h3F1E, 16'h001E,
16'h3F1F, 16'h001F



};


endpackage
