


module nametable_decoder_tb();

reg [8:0] screen_pixel_row, screen_pixel_col;

reg [15:0] cpu_scroll_addr;




initial begin




end




endmodule